magic
tech sky130A
magscale 1 2
timestamp 1736083967
<< nwell >>
rect -466 -1862 466 1862
<< mvpmos >>
rect -208 -1564 -108 1636
rect -50 -1564 50 1636
rect 108 -1564 208 1636
<< mvpdiff >>
rect -266 1624 -208 1636
rect -266 -1552 -254 1624
rect -220 -1552 -208 1624
rect -266 -1564 -208 -1552
rect -108 1624 -50 1636
rect -108 -1552 -96 1624
rect -62 -1552 -50 1624
rect -108 -1564 -50 -1552
rect 50 1624 108 1636
rect 50 -1552 62 1624
rect 96 -1552 108 1624
rect 50 -1564 108 -1552
rect 208 1624 266 1636
rect 208 -1552 220 1624
rect 254 -1552 266 1624
rect 208 -1564 266 -1552
<< mvpdiffc >>
rect -254 -1552 -220 1624
rect -96 -1552 -62 1624
rect 62 -1552 96 1624
rect 220 -1552 254 1624
<< mvnsubdiff >>
rect -400 1784 400 1796
rect -400 1750 -292 1784
rect 292 1750 400 1784
rect -400 1738 400 1750
rect -400 -1738 -342 1738
rect 342 -1738 400 1738
rect -400 -1750 400 -1738
rect -400 -1784 -292 -1750
rect 292 -1784 400 -1750
rect -400 -1796 400 -1784
<< mvnsubdiffcont >>
rect -292 1750 292 1784
rect -292 -1784 292 -1750
<< poly >>
rect -208 1636 -108 1662
rect -50 1636 50 1662
rect 108 1636 208 1662
rect -208 -1611 -108 -1564
rect -208 -1645 -192 -1611
rect -124 -1645 -108 -1611
rect -208 -1661 -108 -1645
rect -50 -1611 50 -1564
rect -50 -1645 -34 -1611
rect 34 -1645 50 -1611
rect -50 -1661 50 -1645
rect 108 -1611 208 -1564
rect 108 -1645 124 -1611
rect 192 -1645 208 -1611
rect 108 -1661 208 -1645
<< polycont >>
rect -192 -1645 -124 -1611
rect -34 -1645 34 -1611
rect 124 -1645 192 -1611
<< locali >>
rect -308 1750 -292 1784
rect 292 1750 308 1784
rect -254 1624 -220 1640
rect -254 -1568 -220 -1552
rect -96 1624 -62 1640
rect -96 -1568 -62 -1552
rect 62 1624 96 1640
rect 62 -1568 96 -1552
rect 220 1624 254 1640
rect 220 -1568 254 -1552
rect -208 -1645 -192 -1611
rect -124 -1645 -108 -1611
rect -50 -1645 -34 -1611
rect 34 -1645 50 -1611
rect 108 -1645 124 -1611
rect 192 -1645 208 -1611
rect -308 -1784 -292 -1750
rect 292 -1784 308 -1750
<< viali >>
rect -254 -1552 -220 1624
rect -96 -1552 -62 1624
rect 62 -1552 96 1624
rect 220 -1552 254 1624
rect -192 -1645 -124 -1611
rect -34 -1645 34 -1611
rect 124 -1645 192 -1611
<< metal1 >>
rect -260 1624 -214 1636
rect -260 -1552 -254 1624
rect -220 -1552 -214 1624
rect -260 -1564 -214 -1552
rect -102 1624 -56 1636
rect -102 -1552 -96 1624
rect -62 -1552 -56 1624
rect -102 -1564 -56 -1552
rect 56 1624 102 1636
rect 56 -1552 62 1624
rect 96 -1552 102 1624
rect 56 -1564 102 -1552
rect 214 1624 260 1636
rect 214 -1552 220 1624
rect 254 -1552 260 1624
rect 214 -1564 260 -1552
rect -204 -1611 -112 -1605
rect -204 -1645 -192 -1611
rect -124 -1645 -112 -1611
rect -204 -1651 -112 -1645
rect -46 -1611 46 -1605
rect -46 -1645 -34 -1611
rect 34 -1645 46 -1611
rect -46 -1651 46 -1645
rect 112 -1611 204 -1605
rect 112 -1645 124 -1611
rect 192 -1645 204 -1611
rect 112 -1651 204 -1645
<< properties >>
string FIXED_BBOX -371 -1767 371 1767
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 16.0 l 0.5 m 1 nf 3 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
