magic
tech sky130A
magscale 1 2
timestamp 1735905388
<< error_p >>
rect -1127 -316 -1097 316
rect -1061 -250 -1031 250
rect 1031 -250 1061 250
rect 1097 -316 1127 316
<< nwell >>
rect -1097 -350 1097 350
<< mvpmos >>
rect -1003 -250 -803 250
rect -745 -250 -545 250
rect -487 -250 -287 250
rect -229 -250 -29 250
rect 29 -250 229 250
rect 287 -250 487 250
rect 545 -250 745 250
rect 803 -250 1003 250
<< mvpdiff >>
rect -1061 238 -1003 250
rect -1061 -238 -1049 238
rect -1015 -238 -1003 238
rect -1061 -250 -1003 -238
rect -803 238 -745 250
rect -803 -238 -791 238
rect -757 -238 -745 238
rect -803 -250 -745 -238
rect -545 238 -487 250
rect -545 -238 -533 238
rect -499 -238 -487 238
rect -545 -250 -487 -238
rect -287 238 -229 250
rect -287 -238 -275 238
rect -241 -238 -229 238
rect -287 -250 -229 -238
rect -29 238 29 250
rect -29 -238 -17 238
rect 17 -238 29 238
rect -29 -250 29 -238
rect 229 238 287 250
rect 229 -238 241 238
rect 275 -238 287 238
rect 229 -250 287 -238
rect 487 238 545 250
rect 487 -238 499 238
rect 533 -238 545 238
rect 487 -250 545 -238
rect 745 238 803 250
rect 745 -238 757 238
rect 791 -238 803 238
rect 745 -250 803 -238
rect 1003 238 1061 250
rect 1003 -238 1015 238
rect 1049 -238 1061 238
rect 1003 -250 1061 -238
<< mvpdiffc >>
rect -1049 -238 -1015 238
rect -791 -238 -757 238
rect -533 -238 -499 238
rect -275 -238 -241 238
rect -17 -238 17 238
rect 241 -238 275 238
rect 499 -238 533 238
rect 757 -238 791 238
rect 1015 -238 1049 238
<< poly >>
rect -1003 331 -803 347
rect -1003 297 -987 331
rect -819 297 -803 331
rect -1003 250 -803 297
rect -745 331 -545 347
rect -745 297 -729 331
rect -561 297 -545 331
rect -745 250 -545 297
rect -487 331 -287 347
rect -487 297 -471 331
rect -303 297 -287 331
rect -487 250 -287 297
rect -229 331 -29 347
rect -229 297 -213 331
rect -45 297 -29 331
rect -229 250 -29 297
rect 29 331 229 347
rect 29 297 45 331
rect 213 297 229 331
rect 29 250 229 297
rect 287 331 487 347
rect 287 297 303 331
rect 471 297 487 331
rect 287 250 487 297
rect 545 331 745 347
rect 545 297 561 331
rect 729 297 745 331
rect 545 250 745 297
rect 803 331 1003 347
rect 803 297 819 331
rect 987 297 1003 331
rect 803 250 1003 297
rect -1003 -297 -803 -250
rect -1003 -331 -987 -297
rect -819 -331 -803 -297
rect -1003 -347 -803 -331
rect -745 -297 -545 -250
rect -745 -331 -729 -297
rect -561 -331 -545 -297
rect -745 -347 -545 -331
rect -487 -297 -287 -250
rect -487 -331 -471 -297
rect -303 -331 -287 -297
rect -487 -347 -287 -331
rect -229 -297 -29 -250
rect -229 -331 -213 -297
rect -45 -331 -29 -297
rect -229 -347 -29 -331
rect 29 -297 229 -250
rect 29 -331 45 -297
rect 213 -331 229 -297
rect 29 -347 229 -331
rect 287 -297 487 -250
rect 287 -331 303 -297
rect 471 -331 487 -297
rect 287 -347 487 -331
rect 545 -297 745 -250
rect 545 -331 561 -297
rect 729 -331 745 -297
rect 545 -347 745 -331
rect 803 -297 1003 -250
rect 803 -331 819 -297
rect 987 -331 1003 -297
rect 803 -347 1003 -331
<< polycont >>
rect -987 297 -819 331
rect -729 297 -561 331
rect -471 297 -303 331
rect -213 297 -45 331
rect 45 297 213 331
rect 303 297 471 331
rect 561 297 729 331
rect 819 297 987 331
rect -987 -331 -819 -297
rect -729 -331 -561 -297
rect -471 -331 -303 -297
rect -213 -331 -45 -297
rect 45 -331 213 -297
rect 303 -331 471 -297
rect 561 -331 729 -297
rect 819 -331 987 -297
<< locali >>
rect -1003 297 -987 331
rect -819 297 -803 331
rect -745 297 -729 331
rect -561 297 -545 331
rect -487 297 -471 331
rect -303 297 -287 331
rect -229 297 -213 331
rect -45 297 -29 331
rect 29 297 45 331
rect 213 297 229 331
rect 287 297 303 331
rect 471 297 487 331
rect 545 297 561 331
rect 729 297 745 331
rect 803 297 819 331
rect 987 297 1003 331
rect -1049 238 -1015 254
rect -1049 -254 -1015 -238
rect -791 238 -757 254
rect -791 -254 -757 -238
rect -533 238 -499 254
rect -533 -254 -499 -238
rect -275 238 -241 254
rect -275 -254 -241 -238
rect -17 238 17 254
rect -17 -254 17 -238
rect 241 238 275 254
rect 241 -254 275 -238
rect 499 238 533 254
rect 499 -254 533 -238
rect 757 238 791 254
rect 757 -254 791 -238
rect 1015 238 1049 254
rect 1015 -254 1049 -238
rect -1003 -331 -987 -297
rect -819 -331 -803 -297
rect -745 -331 -729 -297
rect -561 -331 -545 -297
rect -487 -331 -471 -297
rect -303 -331 -287 -297
rect -229 -331 -213 -297
rect -45 -331 -29 -297
rect 29 -331 45 -297
rect 213 -331 229 -297
rect 287 -331 303 -297
rect 471 -331 487 -297
rect 545 -331 561 -297
rect 729 -331 745 -297
rect 803 -331 819 -297
rect 987 -331 1003 -297
<< viali >>
rect -987 297 -819 331
rect -729 297 -561 331
rect -471 297 -303 331
rect -213 297 -45 331
rect 45 297 213 331
rect 303 297 471 331
rect 561 297 729 331
rect 819 297 987 331
rect -1049 -238 -1015 238
rect -791 -238 -757 238
rect -533 -238 -499 238
rect -275 -238 -241 238
rect -17 -238 17 238
rect 241 -238 275 238
rect 499 -238 533 238
rect 757 -238 791 238
rect 1015 -238 1049 238
rect -987 -331 -819 -297
rect -729 -331 -561 -297
rect -471 -331 -303 -297
rect -213 -331 -45 -297
rect 45 -331 213 -297
rect 303 -331 471 -297
rect 561 -331 729 -297
rect 819 -331 987 -297
<< metal1 >>
rect -999 331 -807 337
rect -999 297 -987 331
rect -819 297 -807 331
rect -999 291 -807 297
rect -741 331 -549 337
rect -741 297 -729 331
rect -561 297 -549 331
rect -741 291 -549 297
rect -483 331 -291 337
rect -483 297 -471 331
rect -303 297 -291 331
rect -483 291 -291 297
rect -225 331 -33 337
rect -225 297 -213 331
rect -45 297 -33 331
rect -225 291 -33 297
rect 33 331 225 337
rect 33 297 45 331
rect 213 297 225 331
rect 33 291 225 297
rect 291 331 483 337
rect 291 297 303 331
rect 471 297 483 331
rect 291 291 483 297
rect 549 331 741 337
rect 549 297 561 331
rect 729 297 741 331
rect 549 291 741 297
rect 807 331 999 337
rect 807 297 819 331
rect 987 297 999 331
rect 807 291 999 297
rect -1055 238 -1009 250
rect -1055 -238 -1049 238
rect -1015 -238 -1009 238
rect -1055 -250 -1009 -238
rect -797 238 -751 250
rect -797 -238 -791 238
rect -757 -238 -751 238
rect -797 -250 -751 -238
rect -539 238 -493 250
rect -539 -238 -533 238
rect -499 -238 -493 238
rect -539 -250 -493 -238
rect -281 238 -235 250
rect -281 -238 -275 238
rect -241 -238 -235 238
rect -281 -250 -235 -238
rect -23 238 23 250
rect -23 -238 -17 238
rect 17 -238 23 238
rect -23 -250 23 -238
rect 235 238 281 250
rect 235 -238 241 238
rect 275 -238 281 238
rect 235 -250 281 -238
rect 493 238 539 250
rect 493 -238 499 238
rect 533 -238 539 238
rect 493 -250 539 -238
rect 751 238 797 250
rect 751 -238 757 238
rect 791 -238 797 238
rect 751 -250 797 -238
rect 1009 238 1055 250
rect 1009 -238 1015 238
rect 1049 -238 1055 238
rect 1009 -250 1055 -238
rect -999 -297 -807 -291
rect -999 -331 -987 -297
rect -819 -331 -807 -297
rect -999 -337 -807 -331
rect -741 -297 -549 -291
rect -741 -331 -729 -297
rect -561 -331 -549 -297
rect -741 -337 -549 -331
rect -483 -297 -291 -291
rect -483 -331 -471 -297
rect -303 -331 -291 -297
rect -483 -337 -291 -331
rect -225 -297 -33 -291
rect -225 -331 -213 -297
rect -45 -331 -33 -297
rect -225 -337 -33 -331
rect 33 -297 225 -291
rect 33 -331 45 -297
rect 213 -331 225 -297
rect 33 -337 225 -331
rect 291 -297 483 -291
rect 291 -331 303 -297
rect 471 -331 483 -297
rect 291 -337 483 -331
rect 549 -297 741 -291
rect 549 -331 561 -297
rect 729 -331 741 -297
rect 549 -337 741 -331
rect 807 -297 999 -291
rect 807 -331 819 -297
rect 987 -331 999 -297
rect 807 -337 999 -331
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 2.5 l 1.0 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
