magic
tech sky130A
magscale 1 2
timestamp 1736115234
<< pwell >>
rect 2332 -2894 2400 -636
rect 2332 -2980 8836 -2894
<< viali >>
rect 2354 -2872 2388 -572
rect 8802 -2872 8836 -572
rect 2450 -2968 8740 -2934
<< metal1 >>
rect 2332 -572 2848 -400
rect 2332 -2872 2354 -572
rect 2388 -1034 2848 -572
rect 3392 -606 3592 -406
rect 4092 -604 4292 -404
rect 4790 -604 4990 -404
rect 5496 -604 5696 -404
rect 6196 -602 6396 -402
rect 6896 -602 7096 -402
rect 7598 -602 7798 -402
rect 2962 -1034 3314 -612
rect 3430 -1034 3548 -606
rect 3666 -1030 4014 -608
rect 2388 -2872 2612 -1034
rect 3194 -2180 3314 -1034
rect 3666 -1036 4018 -1030
rect 4128 -1036 4252 -604
rect 4368 -1036 4726 -612
rect 4830 -1030 4952 -604
rect 5066 -1032 5420 -608
rect 3194 -2300 3782 -2180
rect 2728 -2832 3080 -2410
rect 3198 -2834 3550 -2412
rect 3660 -2556 3782 -2300
rect 3900 -2186 4018 -1036
rect 4598 -2172 4726 -1036
rect 3900 -2191 4487 -2186
rect 3900 -2304 4488 -2191
rect 4598 -2300 5192 -2172
rect 5300 -2180 5420 -1032
rect 5536 -1034 5656 -604
rect 5772 -1034 6122 -612
rect 6238 -1034 6356 -602
rect 6470 -612 6822 -610
rect 6470 -1034 6824 -612
rect 6940 -1034 7058 -602
rect 7170 -1034 7526 -610
rect 7642 -1034 7760 -602
rect 7876 -1034 8228 -400
rect 8302 -602 8502 -402
rect 8578 -572 8858 -440
rect 8344 -1034 8462 -602
rect 6000 -2180 6122 -1034
rect 6700 -2180 6824 -1034
rect 7400 -2174 7526 -1034
rect 5300 -2300 5888 -2180
rect 3660 -2564 3780 -2556
rect 3660 -2832 3722 -2564
rect 3894 -2838 4250 -2408
rect 4366 -2832 4488 -2304
rect 4598 -2834 4956 -2410
rect 5064 -2832 5192 -2300
rect 5302 -2834 5656 -2410
rect 5766 -2832 5888 -2300
rect 6000 -2302 6592 -2180
rect 6700 -2300 7294 -2180
rect 7400 -2246 7999 -2174
rect 7400 -2300 8000 -2246
rect 6004 -2832 6354 -2410
rect 6468 -2832 6592 -2302
rect 6706 -2832 7060 -2410
rect 7172 -2832 7294 -2300
rect 7408 -2832 7760 -2412
rect 7870 -2832 8000 -2300
rect 8110 -2832 8462 -2410
rect 2332 -2888 2612 -2872
rect 8578 -2872 8802 -572
rect 8836 -2872 8858 -572
rect 8578 -2888 8858 -2872
rect 2332 -2934 8858 -2888
rect 2332 -2968 2450 -2934
rect 8740 -2968 8858 -2934
rect 2332 -2980 8858 -2968
use sky130_fd_pr__res_xhigh_po_0p69_C3M8XK  XR1
timestamp 1736113453
transform 1 0 5595 0 1 -1722
box -3277 -1282 3277 1282
<< labels >>
flabel metal1 2332 -600 2532 -400 0 FreeSans 256 0 0 0 COM
port 8 nsew
flabel metal1 7956 -600 8156 -400 0 FreeSans 256 0 0 0 OUT
port 9 nsew
flabel metal1 3392 -606 3592 -406 0 FreeSans 256 0 0 0 B0
port 1 nsew
flabel metal1 4092 -604 4292 -404 0 FreeSans 256 0 0 0 B1
port 0 nsew
flabel metal1 4790 -604 4990 -404 0 FreeSans 256 0 0 0 B2
port 2 nsew
flabel metal1 5496 -604 5696 -404 0 FreeSans 256 0 0 0 B3
port 3 nsew
flabel metal1 6196 -602 6396 -402 0 FreeSans 256 0 0 0 B4
port 5 nsew
flabel metal1 6896 -602 7096 -402 0 FreeSans 256 0 0 0 B5
port 7 nsew
flabel metal1 7598 -602 7798 -402 0 FreeSans 256 0 0 0 B6
port 6 nsew
flabel metal1 8302 -602 8502 -402 0 FreeSans 256 0 0 0 B7
port 4 nsew
<< end >>
