magic
tech sky130A
magscale 1 2
timestamp 1736799799
<< mvnmos >>
rect -629 -100 -29 100
rect 29 -100 629 100
<< mvndiff >>
rect -687 88 -629 100
rect -687 -88 -675 88
rect -641 -88 -629 88
rect -687 -100 -629 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 629 88 687 100
rect 629 -88 641 88
rect 675 -88 687 88
rect 629 -100 687 -88
<< mvndiffc >>
rect -675 -88 -641 88
rect -17 -88 17 88
rect 641 -88 675 88
<< poly >>
rect -629 172 -29 188
rect -629 138 -613 172
rect -45 138 -29 172
rect -629 100 -29 138
rect 29 172 629 188
rect 29 138 45 172
rect 613 138 629 172
rect 29 100 629 138
rect -629 -138 -29 -100
rect -629 -172 -613 -138
rect -45 -172 -29 -138
rect -629 -188 -29 -172
rect 29 -138 629 -100
rect 29 -172 45 -138
rect 613 -172 629 -138
rect 29 -188 629 -172
<< polycont >>
rect -613 138 -45 172
rect 45 138 613 172
rect -613 -172 -45 -138
rect 45 -172 613 -138
<< locali >>
rect -629 138 -613 172
rect -45 138 -29 172
rect 29 138 45 172
rect 613 138 629 172
rect -675 88 -641 104
rect -675 -104 -641 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 641 88 675 104
rect 641 -104 675 -88
rect -629 -172 -613 -138
rect -45 -172 -29 -138
rect 29 -172 45 -138
rect 613 -172 629 -138
<< viali >>
rect -613 138 -45 172
rect 45 138 613 172
rect -675 -88 -641 88
rect -17 -88 17 88
rect 641 -88 675 88
rect -613 -172 -45 -138
rect 45 -172 613 -138
<< metal1 >>
rect -625 172 -33 178
rect -625 138 -613 172
rect -45 138 -33 172
rect -625 132 -33 138
rect 33 172 625 178
rect 33 138 45 172
rect 613 138 625 172
rect 33 132 625 138
rect -681 88 -635 100
rect -681 -88 -675 88
rect -641 -88 -635 88
rect -681 -100 -635 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 635 88 681 100
rect 635 -88 641 88
rect 675 -88 681 88
rect 635 -100 681 -88
rect -625 -138 -33 -132
rect -625 -172 -613 -138
rect -45 -172 -33 -138
rect -625 -178 -33 -172
rect 33 -138 625 -132
rect 33 -172 45 -138
rect 613 -172 625 -138
rect 33 -178 625 -172
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 3.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
