magic
tech sky130A
magscale 1 2
timestamp 1736094482
<< pwell >>
rect 1106 -1246 1152 -1108
rect 1106 -1260 1150 -1246
<< locali >>
rect 1016 274 1400 308
<< viali >>
rect 900 4222 1516 4256
rect 900 -1312 1516 -1278
<< metal1 >>
rect 808 4256 1608 4390
rect 808 4222 900 4256
rect 1516 4222 1608 4256
rect 808 4190 1608 4222
rect 948 908 994 4190
rect 1090 908 1100 4110
rect 1158 908 1168 4110
rect 1264 908 1310 4190
rect 1406 908 1416 4108
rect 1474 908 1484 4108
rect 1004 668 1096 868
rect 1162 668 1254 868
rect 1320 668 1412 868
rect 1004 468 1412 668
rect 1004 268 1096 468
rect 1162 268 1254 468
rect 1320 268 1412 468
rect 1090 -1164 1100 236
rect 1158 -1164 1168 236
rect 1406 -1164 1416 236
rect 1474 -1164 1484 236
rect 948 -1246 994 -1164
rect 1264 -1246 1310 -1164
rect 808 -1278 1608 -1246
rect 808 -1312 900 -1278
rect 1516 -1312 1608 -1278
rect 808 -1446 1608 -1312
<< via1 >>
rect 1100 908 1158 4110
rect 1416 908 1474 4108
rect 1100 -1164 1158 236
rect 1416 -1164 1474 236
<< metal2 >>
rect 1100 4110 1158 4120
rect 1100 236 1158 908
rect 1100 -1246 1158 -1164
rect 1416 4108 1474 4118
rect 1416 236 1474 908
rect 1416 -1246 1474 -1164
rect 1100 -1446 1474 -1246
use sky130_fd_pr__pfet_g5v0d10v5_U8PLV5  sky130_fd_pr__pfet_g5v0d10v5_U8PLV5_0
timestamp 1736083967
transform 1 0 1208 0 1 2472
box -466 -1862 466 1862
use sky130_fd_pr__nfet_g5v0d10v5_GUT4ZJ  XM2
timestamp 1736083967
transform 1 0 1208 0 1 -433
box -436 -927 436 927
<< labels >>
flabel metal1 1108 468 1308 668 0 FreeSans 256 0 0 0 Dx
port 1 nsew
flabel metal1 808 4190 1008 4390 0 FreeSans 256 0 0 0 Vref
port 0 nsew
flabel metal1 808 -1446 1008 -1246 0 FreeSans 256 0 0 0 Vcom
port 3 nsew
flabel metal2 1190 -1446 1390 -1246 0 FreeSans 256 0 0 0 Outx
port 2 nsew
<< end >>
