magic
tech sky130A
magscale 1 2
timestamp 1735905531
<< error_p >>
rect -353 -2566 -323 2566
rect -287 -2500 -257 2500
rect 257 -2500 287 2500
rect 323 -2566 353 2566
<< nwell >>
rect -323 -2600 323 2600
<< mvpmos >>
rect -229 -2500 -29 2500
rect 29 -2500 229 2500
<< mvpdiff >>
rect -287 2488 -229 2500
rect -287 -2488 -275 2488
rect -241 -2488 -229 2488
rect -287 -2500 -229 -2488
rect -29 2488 29 2500
rect -29 -2488 -17 2488
rect 17 -2488 29 2488
rect -29 -2500 29 -2488
rect 229 2488 287 2500
rect 229 -2488 241 2488
rect 275 -2488 287 2488
rect 229 -2500 287 -2488
<< mvpdiffc >>
rect -275 -2488 -241 2488
rect -17 -2488 17 2488
rect 241 -2488 275 2488
<< poly >>
rect -229 2581 -29 2597
rect -229 2547 -213 2581
rect -45 2547 -29 2581
rect -229 2500 -29 2547
rect 29 2581 229 2597
rect 29 2547 45 2581
rect 213 2547 229 2581
rect 29 2500 229 2547
rect -229 -2547 -29 -2500
rect -229 -2581 -213 -2547
rect -45 -2581 -29 -2547
rect -229 -2597 -29 -2581
rect 29 -2547 229 -2500
rect 29 -2581 45 -2547
rect 213 -2581 229 -2547
rect 29 -2597 229 -2581
<< polycont >>
rect -213 2547 -45 2581
rect 45 2547 213 2581
rect -213 -2581 -45 -2547
rect 45 -2581 213 -2547
<< locali >>
rect -229 2547 -213 2581
rect -45 2547 -29 2581
rect 29 2547 45 2581
rect 213 2547 229 2581
rect -275 2488 -241 2504
rect -275 -2504 -241 -2488
rect -17 2488 17 2504
rect -17 -2504 17 -2488
rect 241 2488 275 2504
rect 241 -2504 275 -2488
rect -229 -2581 -213 -2547
rect -45 -2581 -29 -2547
rect 29 -2581 45 -2547
rect 213 -2581 229 -2547
<< viali >>
rect -213 2547 -45 2581
rect 45 2547 213 2581
rect -275 -2488 -241 2488
rect -17 -2488 17 2488
rect 241 -2488 275 2488
rect -213 -2581 -45 -2547
rect 45 -2581 213 -2547
<< metal1 >>
rect -225 2581 -33 2587
rect -225 2547 -213 2581
rect -45 2547 -33 2581
rect -225 2541 -33 2547
rect 33 2581 225 2587
rect 33 2547 45 2581
rect 213 2547 225 2581
rect 33 2541 225 2547
rect -281 2488 -235 2500
rect -281 -2488 -275 2488
rect -241 -2488 -235 2488
rect -281 -2500 -235 -2488
rect -23 2488 23 2500
rect -23 -2488 -17 2488
rect 17 -2488 23 2488
rect -23 -2500 23 -2488
rect 235 2488 281 2500
rect 235 -2488 241 2488
rect 275 -2488 281 2488
rect 235 -2500 281 -2488
rect -225 -2547 -33 -2541
rect -225 -2581 -213 -2547
rect -45 -2581 -33 -2547
rect -225 -2587 -33 -2581
rect 33 -2547 225 -2541
rect 33 -2581 45 -2547
rect 213 -2581 225 -2547
rect 33 -2587 225 -2581
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 25.0 l 1.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
