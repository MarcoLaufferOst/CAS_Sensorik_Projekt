magic
tech sky130A
magscale 1 2
timestamp 1737189919
<< nwell >>
rect 940 3830 16070 4710
rect 940 2830 13680 3830
<< mvpsubdiff >>
rect 16160 4620 23570 4640
rect 16160 4540 16260 4620
rect 23360 4540 23570 4620
rect 16160 4520 23570 4540
rect 16160 3740 16280 4520
rect 13770 3620 16280 3740
rect 13770 2890 13890 3620
rect 23450 2890 23570 4520
rect 13770 2870 23570 2890
rect 13770 2790 13870 2870
rect 23380 2790 23570 2870
rect 13770 2770 23570 2790
rect 1010 1850 23780 1870
rect 1010 1770 1110 1850
rect 23680 1770 23780 1850
rect 1010 1750 23780 1770
rect 1010 -540 1130 1750
rect 23660 -540 23780 1750
rect 1010 -560 23780 -540
rect 1010 -640 1110 -560
rect 23680 -640 23780 -560
rect 1010 -660 23780 -640
<< mvnsubdiff >>
rect 1010 4620 15970 4640
rect 1010 4540 1110 4620
rect 15870 4540 15970 4620
rect 1010 4520 15970 4540
rect 1010 3020 1130 4520
rect 13490 4040 13610 4520
rect 15850 4040 15970 4520
rect 13490 3920 15970 4040
rect 13490 3020 13610 3920
rect 1010 3000 13610 3020
rect 1010 2920 1110 3000
rect 13510 2920 13610 3000
rect 1010 2900 13610 2920
<< mvpsubdiffcont >>
rect 16260 4540 23360 4620
rect 13870 2790 23380 2870
rect 1110 1770 23680 1850
rect 1110 -640 23680 -560
<< mvnsubdiffcont >>
rect 1110 4540 15870 4620
rect 1110 2920 13510 3000
<< locali >>
rect 1030 2920 1110 4620
rect 13510 4020 13590 4540
rect 15870 4020 15950 4620
rect 13510 3940 15950 4020
rect 13510 2920 13590 3940
rect 16180 3720 16260 4620
rect 23360 4540 23550 4620
rect 13790 3640 16260 3720
rect 13790 2790 13870 3640
rect 23470 2870 23550 4540
rect 23380 2790 23550 2870
rect 1030 -640 1110 1850
rect 23680 -640 23760 1850
<< viali >>
rect 1110 4540 15870 4620
rect 1110 2920 13510 3000
rect 16260 4540 23360 4620
rect 13870 2790 23380 2870
rect 1110 1770 23680 1850
rect 1110 -640 23680 -560
<< metal1 >>
rect 940 4810 23570 5080
rect 940 4710 1310 4810
rect 1410 4800 4066 4810
rect 1410 4710 2138 4800
rect 2238 4710 4066 4800
rect 4166 4710 5994 4810
rect 6094 4710 7922 4810
rect 8022 4710 9850 4810
rect 9950 4710 11778 4810
rect 11878 4710 13200 4810
rect 13300 4710 13660 4810
rect 13760 4710 23570 4810
rect 940 4680 23570 4710
rect 1010 4640 1860 4680
rect 1010 4620 15970 4640
rect 1010 4540 1110 4620
rect 15870 4540 15970 4620
rect 1010 4520 15970 4540
rect 1010 3020 1130 4520
rect 1300 4402 1310 4460
rect 1410 4402 1420 4460
rect 2128 4402 2138 4460
rect 2238 4402 2248 4460
rect 4056 4402 4066 4460
rect 4166 4402 4176 4460
rect 5984 4402 5994 4460
rect 6094 4402 6104 4460
rect 7912 4402 7922 4460
rect 8022 4402 8032 4460
rect 9840 4402 9850 4460
rect 9950 4402 9960 4460
rect 11768 4402 11778 4460
rect 11878 4402 11888 4460
rect 13190 4402 13200 4461
rect 13300 4402 13310 4461
rect 1160 4020 1170 4120
rect 1230 4020 1240 4120
rect 13370 4060 13380 4160
rect 13450 4060 13460 4160
rect 13490 4040 13610 4520
rect 13910 4410 13920 4470
rect 14020 4410 14030 4470
rect 13660 4180 13670 4360
rect 13730 4180 13740 4360
rect 15730 4180 15740 4360
rect 15800 4180 15810 4360
rect 13910 4070 13920 4130
rect 14020 4070 14030 4130
rect 15850 4040 15970 4520
rect 13490 3920 15970 4040
rect 16160 4620 23570 4640
rect 16160 4540 16260 4620
rect 23360 4540 23570 4620
rect 16160 4520 23570 4540
rect 1300 3744 1310 3802
rect 1410 3744 1420 3802
rect 2728 3744 2738 3802
rect 2838 3744 2848 3802
rect 4656 3744 4666 3802
rect 4766 3744 4776 3802
rect 6584 3744 6594 3802
rect 6694 3744 6704 3802
rect 8512 3744 8522 3802
rect 8622 3744 8632 3802
rect 10440 3744 10450 3802
rect 10550 3744 10560 3802
rect 12368 3744 12378 3802
rect 12478 3744 12488 3802
rect 13190 3744 13200 3803
rect 13300 3744 13310 3803
rect 1160 3400 1170 3500
rect 1230 3400 1240 3500
rect 13370 3400 13380 3500
rect 13450 3400 13460 3500
rect 1300 3086 1310 3144
rect 1410 3086 1420 3144
rect 2128 3086 2138 3144
rect 2238 3086 2248 3144
rect 4056 3086 4066 3144
rect 4166 3086 4176 3144
rect 5984 3086 5994 3144
rect 6094 3086 6104 3144
rect 7912 3086 7922 3144
rect 8022 3086 8032 3144
rect 9840 3086 9850 3144
rect 9950 3086 9960 3144
rect 11768 3086 11778 3144
rect 11878 3086 11888 3144
rect 13190 3085 13200 3144
rect 13300 3085 13310 3144
rect 13490 3020 13610 3920
rect 16160 3740 16280 4520
rect 16970 4386 16980 4444
rect 17080 4386 17090 4444
rect 17368 4386 17378 4444
rect 17478 4386 17488 4444
rect 18078 4386 18088 4444
rect 18188 4386 18198 4444
rect 18788 4386 18798 4444
rect 18898 4386 18908 4444
rect 19498 4386 19508 4444
rect 19608 4386 19618 4444
rect 20120 4386 20130 4444
rect 20230 4386 20240 4444
rect 20610 4220 20620 4320
rect 20720 4220 20730 4320
rect 23080 4230 23090 4330
rect 23190 4230 23200 4330
rect 16790 4020 16800 4120
rect 16900 4020 16910 4120
rect 20290 4030 20300 4130
rect 20390 4030 20400 4130
rect 1010 3000 13610 3020
rect 1010 2920 1110 3000
rect 13510 2920 13610 3000
rect 1010 2900 13610 2920
rect 13770 3620 16280 3740
rect 16360 3730 16370 3830
rect 16430 3730 16440 3830
rect 16610 3770 16620 4000
rect 16720 3770 16730 4000
rect 20610 3850 20620 3950
rect 20720 3850 20730 3950
rect 23080 3840 23090 3940
rect 23190 3840 23200 3940
rect 16970 3728 16980 3786
rect 17080 3728 17090 3786
rect 17568 3728 17578 3786
rect 17678 3728 17688 3786
rect 18278 3728 18288 3786
rect 18388 3728 18398 3786
rect 18988 3728 18998 3786
rect 19098 3728 19108 3786
rect 19697 3728 19707 3786
rect 19807 3728 19817 3786
rect 20120 3728 20130 3786
rect 20230 3728 20240 3786
rect 13770 2890 13890 3620
rect 14150 3490 14160 3550
rect 14260 3490 14270 3550
rect 13920 3320 13930 3460
rect 14000 3320 14010 3460
rect 16790 3370 16800 3470
rect 16900 3370 16910 3470
rect 20290 3380 20300 3480
rect 20390 3380 20400 3480
rect 20610 3470 20620 3570
rect 20720 3470 20730 3570
rect 23080 3470 23090 3570
rect 23190 3470 23200 3570
rect 15710 3230 15720 3290
rect 15820 3230 15830 3290
rect 16450 3260 16460 3360
rect 16560 3260 16570 3360
rect 13920 3060 13930 3200
rect 14000 3060 14010 3200
rect 16970 3070 16980 3128
rect 17080 3070 17090 3128
rect 17368 3070 17378 3128
rect 17478 3070 17488 3128
rect 18078 3070 18088 3128
rect 18188 3070 18198 3128
rect 18788 3070 18798 3128
rect 18898 3070 18908 3128
rect 19498 3070 19508 3128
rect 19608 3070 19618 3128
rect 20120 3070 20130 3128
rect 20230 3070 20240 3128
rect 20610 3090 20620 3190
rect 20720 3090 20730 3190
rect 23080 3090 23090 3190
rect 23190 3090 23200 3190
rect 14150 2970 14160 3030
rect 14260 2970 14270 3030
rect 23450 2890 23570 4520
rect 13770 2870 23570 2890
rect 13770 2790 13870 2870
rect 23380 2790 23570 2870
rect 13770 2770 23570 2790
rect 13770 2730 13970 2770
rect 940 2630 14160 2730
rect 14260 2630 16620 2730
rect 16720 2630 16980 2730
rect 17080 2630 17378 2730
rect 17478 2630 18088 2730
rect 18188 2630 18798 2730
rect 18898 2630 19508 2730
rect 19608 2630 20130 2730
rect 20230 2630 20620 2730
rect 20720 2630 23570 2730
rect 940 2430 23570 2630
rect 940 2330 1310 2430
rect 1410 2330 11800 2430
rect 11900 2330 23390 2430
rect 23490 2330 23570 2430
rect 1370 1870 1570 2330
rect 1010 1850 23780 1870
rect 1010 1770 1110 1850
rect 23680 1770 23780 1850
rect 1010 1750 23780 1770
rect 1010 -540 1130 1750
rect 1300 1604 1310 1662
rect 1410 1604 1420 1662
rect 2460 1604 2470 1662
rect 2570 1604 2580 1662
rect 5570 1604 5580 1662
rect 5680 1604 5690 1662
rect 8680 1604 8690 1662
rect 8790 1604 8800 1662
rect 11790 1604 11800 1662
rect 11900 1604 11910 1662
rect 14900 1604 14910 1662
rect 15010 1604 15020 1662
rect 18010 1604 18020 1662
rect 18120 1604 18130 1662
rect 21120 1604 21130 1662
rect 21230 1604 21240 1662
rect 23380 1604 23390 1662
rect 23490 1604 23500 1662
rect 1160 1430 1170 1570
rect 1240 1430 1250 1570
rect 23540 1430 23550 1570
rect 23620 1430 23630 1570
rect 1300 1346 1310 1404
rect 1410 1346 1420 1404
rect 3460 1346 3470 1404
rect 3570 1346 3580 1404
rect 6570 1346 6580 1404
rect 6680 1346 6690 1404
rect 9680 1346 9690 1404
rect 9790 1346 9800 1404
rect 12790 1346 12800 1404
rect 12900 1346 12910 1404
rect 15900 1346 15910 1404
rect 16010 1346 16020 1404
rect 19010 1346 19020 1404
rect 19120 1346 19130 1404
rect 22120 1346 22130 1404
rect 22230 1346 22240 1404
rect 23380 1346 23390 1404
rect 23490 1346 23500 1404
rect 1160 1180 1170 1320
rect 1240 1180 1250 1320
rect 23540 1180 23550 1320
rect 23620 1180 23630 1320
rect 1300 1088 1310 1146
rect 1410 1088 1420 1146
rect 2460 1088 2470 1146
rect 2570 1088 2580 1146
rect 5570 1088 5580 1146
rect 5680 1088 5690 1146
rect 8680 1088 8690 1146
rect 8790 1088 8800 1146
rect 11790 1088 11800 1146
rect 11900 1088 11910 1146
rect 14900 1088 14910 1146
rect 15010 1088 15020 1146
rect 18010 1088 18020 1146
rect 18120 1088 18130 1146
rect 21120 1088 21130 1146
rect 21230 1088 21240 1146
rect 23380 1088 23390 1146
rect 23490 1088 23500 1146
rect 1160 920 1170 1060
rect 1240 920 1250 1060
rect 23540 920 23550 1060
rect 23620 920 23630 1060
rect 1300 830 1310 888
rect 1410 830 1420 888
rect 3460 830 3470 888
rect 3570 830 3580 888
rect 6570 830 6580 888
rect 6680 830 6690 888
rect 9680 830 9690 888
rect 9790 830 9800 888
rect 12790 830 12800 888
rect 12900 830 12910 888
rect 15900 830 15910 888
rect 16010 830 16020 888
rect 19010 830 19020 888
rect 19120 830 19130 888
rect 22120 830 22130 888
rect 22230 830 22240 888
rect 23380 830 23390 888
rect 23490 830 23500 888
rect 1160 660 1170 800
rect 1240 660 1250 800
rect 23540 660 23550 800
rect 23620 660 23630 800
rect 1300 572 1310 630
rect 1410 572 1420 630
rect 2460 572 2470 630
rect 2570 572 2580 630
rect 5570 572 5580 630
rect 5680 572 5690 630
rect 8680 572 8690 630
rect 8790 572 8800 630
rect 11790 572 11800 630
rect 11900 572 11910 630
rect 14900 572 14910 630
rect 15010 572 15020 630
rect 18010 572 18020 630
rect 18120 572 18130 630
rect 21120 572 21130 630
rect 21230 572 21240 630
rect 23380 572 23390 630
rect 23490 572 23500 630
rect 1160 400 1170 540
rect 1240 400 1250 540
rect 23540 410 23550 550
rect 23620 410 23630 550
rect 1300 314 1310 372
rect 1410 314 1420 372
rect 3460 314 3470 372
rect 3570 314 3580 372
rect 6570 314 6580 372
rect 6680 314 6690 372
rect 9680 314 9690 372
rect 9790 314 9800 372
rect 12790 314 12800 372
rect 12900 314 12910 372
rect 15900 314 15910 372
rect 16010 314 16020 372
rect 19010 314 19020 372
rect 19120 314 19130 372
rect 22120 314 22130 372
rect 22230 314 22240 372
rect 23380 314 23390 372
rect 23490 314 23500 372
rect 1160 140 1170 280
rect 1240 140 1250 280
rect 23540 150 23550 290
rect 23620 150 23630 290
rect 1300 56 1310 114
rect 1410 56 1420 114
rect 2460 56 2470 114
rect 2570 56 2580 114
rect 5570 56 5580 114
rect 5680 56 5690 114
rect 8680 56 8690 114
rect 8790 56 8800 114
rect 11790 56 11800 114
rect 11900 56 11910 114
rect 14900 56 14910 114
rect 15010 56 15020 114
rect 18010 56 18020 114
rect 18120 56 18130 114
rect 21120 56 21130 114
rect 21230 56 21240 114
rect 23380 56 23390 114
rect 23490 56 23500 114
rect 1160 -110 1170 30
rect 1240 -110 1250 30
rect 23540 -110 23550 30
rect 23620 -110 23630 30
rect 1300 -202 1310 -144
rect 1410 -202 1420 -144
rect 3460 -202 3470 -144
rect 3570 -202 3580 -144
rect 6570 -202 6580 -144
rect 6680 -202 6690 -144
rect 9680 -202 9690 -144
rect 9790 -202 9800 -144
rect 12790 -202 12800 -144
rect 12900 -202 12910 -144
rect 15900 -202 15910 -144
rect 16010 -202 16020 -144
rect 19010 -202 19020 -144
rect 19120 -202 19130 -144
rect 22120 -202 22130 -144
rect 22230 -202 22240 -144
rect 23380 -202 23390 -144
rect 23490 -202 23500 -144
rect 1160 -370 1170 -230
rect 1240 -370 1250 -230
rect 23540 -370 23550 -230
rect 23620 -370 23630 -230
rect 1300 -460 1310 -403
rect 1410 -460 1420 -403
rect 2460 -460 2470 -402
rect 2570 -460 2580 -402
rect 5570 -460 5580 -402
rect 5680 -460 5690 -402
rect 8680 -460 8690 -402
rect 8790 -460 8800 -402
rect 11790 -460 11800 -402
rect 11900 -460 11910 -402
rect 14900 -460 14910 -402
rect 15010 -460 15020 -402
rect 18010 -460 18020 -402
rect 18120 -460 18130 -402
rect 21120 -460 21130 -402
rect 21230 -460 21240 -402
rect 23380 -460 23390 -402
rect 23490 -460 23500 -402
rect 23660 -540 23780 1750
rect 1010 -560 23780 -540
rect 1010 -640 1110 -560
rect 23680 -640 23780 -560
rect 1010 -660 23780 -640
<< via1 >>
rect 1310 4710 1410 4810
rect 2138 4710 2238 4800
rect 4066 4710 4166 4810
rect 5994 4710 6094 4810
rect 7922 4710 8022 4810
rect 9850 4710 9950 4810
rect 11778 4710 11878 4810
rect 13200 4710 13300 4810
rect 13660 4710 13760 4810
rect 1310 4402 1410 4460
rect 2138 4402 2238 4460
rect 4066 4402 4166 4460
rect 5994 4402 6094 4460
rect 7922 4402 8022 4460
rect 9850 4402 9950 4460
rect 11778 4402 11878 4460
rect 13200 4402 13300 4461
rect 1170 4020 1230 4120
rect 13380 4060 13450 4160
rect 13920 4410 14020 4470
rect 13670 4180 13730 4360
rect 15740 4180 15800 4360
rect 13920 4070 14020 4130
rect 1310 3744 1410 3802
rect 2738 3744 2838 3802
rect 4666 3744 4766 3802
rect 6594 3744 6694 3802
rect 8522 3744 8622 3802
rect 10450 3744 10550 3802
rect 12378 3744 12478 3802
rect 13200 3744 13300 3803
rect 1170 3400 1230 3500
rect 13380 3400 13450 3500
rect 1310 3086 1410 3144
rect 2138 3086 2238 3144
rect 4066 3086 4166 3144
rect 5994 3086 6094 3144
rect 7922 3086 8022 3144
rect 9850 3086 9950 3144
rect 11778 3086 11878 3144
rect 13200 3085 13300 3144
rect 16980 4386 17080 4444
rect 17378 4386 17478 4444
rect 18088 4386 18188 4444
rect 18798 4386 18898 4444
rect 19508 4386 19608 4444
rect 20130 4386 20230 4444
rect 20620 4220 20720 4320
rect 23090 4230 23190 4330
rect 16800 4020 16900 4120
rect 20300 4030 20390 4130
rect 16370 3730 16430 3830
rect 16620 3770 16720 4000
rect 20620 3850 20720 3950
rect 23090 3840 23190 3940
rect 16980 3728 17080 3786
rect 17578 3728 17678 3786
rect 18288 3728 18388 3786
rect 18998 3728 19098 3786
rect 19707 3728 19807 3786
rect 20130 3728 20230 3786
rect 14160 3490 14260 3550
rect 13930 3320 14000 3460
rect 16800 3370 16900 3470
rect 20300 3380 20390 3480
rect 20620 3470 20720 3570
rect 23090 3470 23190 3570
rect 15720 3230 15820 3290
rect 16460 3260 16560 3360
rect 13930 3060 14000 3200
rect 16980 3070 17080 3128
rect 17378 3070 17478 3128
rect 18088 3070 18188 3128
rect 18798 3070 18898 3128
rect 19508 3070 19608 3128
rect 20130 3070 20230 3128
rect 20620 3090 20720 3190
rect 23090 3090 23190 3190
rect 14160 2970 14260 3030
rect 14160 2630 14260 2730
rect 16620 2630 16720 2730
rect 16980 2630 17080 2730
rect 17378 2630 17478 2730
rect 18088 2630 18188 2730
rect 18798 2630 18898 2730
rect 19508 2630 19608 2730
rect 20130 2630 20230 2730
rect 20620 2630 20720 2730
rect 1310 2330 1410 2430
rect 11800 2330 11900 2430
rect 23390 2330 23490 2430
rect 1310 1604 1410 1662
rect 2470 1604 2570 1662
rect 5580 1604 5680 1662
rect 8690 1604 8790 1662
rect 11800 1604 11900 1662
rect 14910 1604 15010 1662
rect 18020 1604 18120 1662
rect 21130 1604 21230 1662
rect 23390 1604 23490 1662
rect 1170 1430 1240 1570
rect 23550 1430 23620 1570
rect 1310 1346 1410 1404
rect 3470 1346 3570 1404
rect 6580 1346 6680 1404
rect 9690 1346 9790 1404
rect 12800 1346 12900 1404
rect 15910 1346 16010 1404
rect 19020 1346 19120 1404
rect 22130 1346 22230 1404
rect 23390 1346 23490 1404
rect 1170 1180 1240 1320
rect 23550 1180 23620 1320
rect 1310 1088 1410 1146
rect 2470 1088 2570 1146
rect 5580 1088 5680 1146
rect 8690 1088 8790 1146
rect 11800 1088 11900 1146
rect 14910 1088 15010 1146
rect 18020 1088 18120 1146
rect 21130 1088 21230 1146
rect 23390 1088 23490 1146
rect 1170 920 1240 1060
rect 23550 920 23620 1060
rect 1310 830 1410 888
rect 3470 830 3570 888
rect 6580 830 6680 888
rect 9690 830 9790 888
rect 12800 830 12900 888
rect 15910 830 16010 888
rect 19020 830 19120 888
rect 22130 830 22230 888
rect 23390 830 23490 888
rect 1170 660 1240 800
rect 23550 660 23620 800
rect 1310 572 1410 630
rect 2470 572 2570 630
rect 5580 572 5680 630
rect 8690 572 8790 630
rect 11800 572 11900 630
rect 14910 572 15010 630
rect 18020 572 18120 630
rect 21130 572 21230 630
rect 23390 572 23490 630
rect 1170 400 1240 540
rect 23550 410 23620 550
rect 1310 314 1410 372
rect 3470 314 3570 372
rect 6580 314 6680 372
rect 9690 314 9790 372
rect 12800 314 12900 372
rect 15910 314 16010 372
rect 19020 314 19120 372
rect 22130 314 22230 372
rect 23390 314 23490 372
rect 1170 140 1240 280
rect 23550 150 23620 290
rect 1310 56 1410 114
rect 2470 56 2570 114
rect 5580 56 5680 114
rect 8690 56 8790 114
rect 11800 56 11900 114
rect 14910 56 15010 114
rect 18020 56 18120 114
rect 21130 56 21230 114
rect 23390 56 23490 114
rect 1170 -110 1240 30
rect 23550 -110 23620 30
rect 1310 -202 1410 -144
rect 3470 -202 3570 -144
rect 6580 -202 6680 -144
rect 9690 -202 9790 -144
rect 12800 -202 12900 -144
rect 15910 -202 16010 -144
rect 19020 -202 19120 -144
rect 22130 -202 22230 -144
rect 23390 -202 23490 -144
rect 1170 -370 1240 -230
rect 23550 -370 23620 -230
rect 1310 -460 1410 -403
rect 2470 -460 2570 -402
rect 5580 -460 5680 -402
rect 8690 -460 8790 -402
rect 11800 -460 11900 -402
rect 14910 -460 15010 -402
rect 18020 -460 18120 -402
rect 21130 -460 21230 -402
rect 23390 -460 23490 -402
<< metal2 >>
rect 1310 4810 1410 4820
rect 4066 4810 4166 4820
rect 1310 4460 1410 4710
rect 1140 4120 1240 4410
rect 1140 4020 1170 4120
rect 1230 4020 1240 4120
rect 1140 3500 1240 4020
rect 1140 3400 1170 3500
rect 1230 3400 1240 3500
rect 940 2570 1040 2580
rect 940 2160 1040 2470
rect 1140 2370 1240 3400
rect 1310 3802 1410 4402
rect 1310 3144 1410 3744
rect 1310 3076 1410 3086
rect 2138 4800 2238 4810
rect 2138 4460 2238 4710
rect 4066 4460 4166 4710
rect 5994 4810 6094 4820
rect 5994 4460 6094 4710
rect 7922 4810 8022 4820
rect 7922 4460 8022 4710
rect 9850 4810 9950 4820
rect 9850 4460 9950 4710
rect 11778 4810 11878 4820
rect 11778 4460 11878 4710
rect 13200 4810 13300 4820
rect 13200 4461 13300 4710
rect 2138 3144 2238 4402
rect 2138 3076 2238 3086
rect 2738 3802 2838 4460
rect 2738 2770 2838 3744
rect 4066 3144 4166 4402
rect 4066 3076 4166 3086
rect 4666 3802 4766 4460
rect 2738 2660 2838 2670
rect 4666 2570 4766 3744
rect 5994 3144 6094 4402
rect 5994 3076 6094 3086
rect 6594 3802 6694 4460
rect 4666 2460 4766 2470
rect 1140 2260 1240 2270
rect 1310 2430 1410 2440
rect 940 2060 1250 2160
rect 1150 1570 1250 2060
rect 1150 1430 1170 1570
rect 1240 1430 1250 1570
rect 1150 1320 1250 1430
rect 1150 1180 1170 1320
rect 1240 1180 1250 1320
rect 1150 1060 1250 1180
rect 1150 920 1170 1060
rect 1240 920 1250 1060
rect 1150 800 1250 920
rect 1150 660 1170 800
rect 1240 660 1250 800
rect 1150 540 1250 660
rect 1150 400 1170 540
rect 1240 400 1250 540
rect 1150 280 1250 400
rect 1150 140 1170 280
rect 1240 140 1250 280
rect 1150 30 1250 140
rect 1150 -110 1170 30
rect 1240 -110 1250 30
rect 1150 -230 1250 -110
rect 1150 -370 1170 -230
rect 1240 -370 1250 -230
rect 1150 -540 1250 -370
rect 1310 1662 1410 2330
rect 3470 2370 3570 2380
rect 1310 1404 1410 1604
rect 1310 1146 1410 1346
rect 1310 888 1410 1088
rect 1310 630 1410 830
rect 1310 372 1410 572
rect 1310 114 1410 314
rect 1310 -144 1410 56
rect 1310 -403 1410 -202
rect 1310 -540 1410 -460
rect 2470 1970 2570 1980
rect 2470 1662 2570 1870
rect 2470 1146 2570 1604
rect 2470 630 2570 1088
rect 2470 114 2570 572
rect 2470 -402 2570 56
rect 2470 -540 2570 -460
rect 3470 1404 3570 2270
rect 6594 2370 6694 3744
rect 7922 3144 8022 4402
rect 7922 3076 8022 3086
rect 8522 3802 8622 4460
rect 6594 2260 6694 2270
rect 6800 2370 6900 2380
rect 6800 2170 6900 2270
rect 8522 2370 8622 3744
rect 9850 3144 9950 4402
rect 9850 3076 9950 3086
rect 10450 3802 10550 4460
rect 10450 2570 10550 3744
rect 11778 3144 11878 4402
rect 11778 3076 11878 3086
rect 12378 3802 12478 4460
rect 12378 2770 12478 3744
rect 13200 3803 13300 4402
rect 13660 4810 13760 4820
rect 13200 3144 13300 3744
rect 13200 3075 13300 3085
rect 13370 4160 13470 4400
rect 13660 4360 13760 4710
rect 13660 4180 13670 4360
rect 13730 4180 13760 4360
rect 13660 4160 13760 4180
rect 13920 4470 14020 4480
rect 13370 4060 13380 4160
rect 13450 4060 13470 4160
rect 13370 3820 13470 4060
rect 13370 3500 13470 3720
rect 13370 3400 13380 3500
rect 13450 3400 13470 3500
rect 13370 2770 13470 3400
rect 12378 2660 12478 2670
rect 13070 2670 13470 2770
rect 13920 4130 14020 4410
rect 16980 4444 17080 4454
rect 13920 3460 14020 4070
rect 15720 4360 15820 4380
rect 15720 4180 15740 4360
rect 15800 4180 15820 4360
rect 13920 3320 13930 3460
rect 14000 3320 14020 3460
rect 13920 3200 14020 3320
rect 13920 3060 13930 3200
rect 14000 3060 14020 3200
rect 10450 2460 10550 2470
rect 12800 2570 12900 2580
rect 11800 2430 11900 2440
rect 8522 2260 8622 2270
rect 9690 2370 9790 2380
rect 6580 2070 6900 2170
rect 3470 888 3570 1346
rect 3470 372 3570 830
rect 3470 -144 3570 314
rect 3470 -540 3570 -202
rect 5580 1970 5680 1980
rect 5580 1662 5680 1870
rect 5580 1146 5680 1604
rect 5580 630 5680 1088
rect 5580 114 5680 572
rect 5580 -402 5680 56
rect 5580 -540 5680 -460
rect 6580 1404 6680 2070
rect 6580 888 6680 1346
rect 6580 372 6680 830
rect 6580 -144 6680 314
rect 6580 -540 6680 -202
rect 8690 1970 8790 1980
rect 8690 1662 8790 1870
rect 8690 1146 8790 1604
rect 8690 630 8790 1088
rect 8690 114 8790 572
rect 8690 -402 8790 56
rect 8690 -540 8790 -460
rect 9690 1404 9790 2270
rect 9690 888 9790 1346
rect 9690 372 9790 830
rect 9690 -144 9790 314
rect 9690 -540 9790 -202
rect 11800 1662 11900 2330
rect 11800 1146 11900 1604
rect 11800 630 11900 1088
rect 11800 114 11900 572
rect 11800 -402 11900 56
rect 11800 -540 11900 -460
rect 12800 1404 12900 2470
rect 13070 2370 13170 2670
rect 13920 2570 14020 3060
rect 14160 3550 14260 3560
rect 14160 3030 14260 3490
rect 15720 3360 15820 4180
rect 16620 4000 16720 4380
rect 16370 3830 16430 3840
rect 16370 3720 16430 3730
rect 16460 3360 16560 3370
rect 16460 3250 16560 3260
rect 15720 2970 15820 3230
rect 14160 2730 14260 2970
rect 14160 2620 14260 2630
rect 16620 2730 16720 3770
rect 16800 4120 16900 4390
rect 16800 3470 16900 4020
rect 16800 2770 16900 3370
rect 16800 2660 16900 2670
rect 16980 3786 17080 4386
rect 16980 3128 17080 3728
rect 16980 2730 17080 3070
rect 16620 2620 16720 2630
rect 16980 2620 17080 2630
rect 17378 4444 17478 4454
rect 17378 3128 17478 4386
rect 17378 2730 17478 3070
rect 17378 2620 17478 2630
rect 17578 3786 17678 4450
rect 13920 2460 14020 2470
rect 13070 2260 13170 2270
rect 15910 2370 16010 2380
rect 12800 888 12900 1346
rect 12800 372 12900 830
rect 12800 -144 12900 314
rect 12800 -540 12900 -202
rect 14910 1970 15010 1980
rect 14910 1662 15010 1870
rect 14910 1146 15010 1604
rect 14910 630 15010 1088
rect 14910 114 15010 572
rect 14910 -402 15010 56
rect 14910 -540 15010 -460
rect 15910 1404 16010 2270
rect 17578 2170 17678 3728
rect 18088 4444 18188 4454
rect 18088 3128 18188 4386
rect 18088 2730 18188 3070
rect 18288 3786 18388 4450
rect 18288 2770 18388 3728
rect 18288 2660 18388 2670
rect 18798 4444 18898 4454
rect 18798 3128 18898 4386
rect 18798 2730 18898 3070
rect 18088 2620 18188 2630
rect 18998 3786 19098 4450
rect 18998 2770 19098 3728
rect 18998 2660 19098 2670
rect 19508 4444 19608 4454
rect 19508 3128 19608 4386
rect 19708 3796 19808 4450
rect 19707 3786 19808 3796
rect 19807 3728 19808 3786
rect 19707 3718 19808 3728
rect 19508 2730 19608 3070
rect 18798 2620 18898 2630
rect 19508 2620 19608 2630
rect 17578 2060 17678 2070
rect 19020 2370 19120 2380
rect 15910 888 16010 1346
rect 15910 372 16010 830
rect 15910 -144 16010 314
rect 15910 -540 16010 -202
rect 18020 1970 18120 1980
rect 18020 1662 18120 1870
rect 18020 1146 18120 1604
rect 18020 630 18120 1088
rect 18020 114 18120 572
rect 18020 -402 18120 56
rect 18020 -540 18120 -460
rect 19020 1404 19120 2270
rect 19708 2170 19808 3718
rect 20130 4444 20230 4454
rect 20130 3786 20230 4386
rect 20130 3128 20230 3728
rect 20130 2730 20230 3070
rect 20290 4130 20390 4390
rect 20290 4030 20300 4130
rect 20290 3480 20390 4030
rect 20290 3380 20300 3480
rect 20290 2770 20390 3380
rect 20290 2660 20390 2670
rect 20620 4320 20720 4420
rect 20620 3950 20720 4220
rect 20620 3570 20720 3850
rect 20620 3190 20720 3470
rect 20620 2730 20720 3090
rect 20130 2620 20230 2630
rect 20620 2620 20720 2630
rect 23090 4330 23190 4420
rect 23090 3940 23190 4230
rect 23090 3570 23190 3840
rect 23090 3190 23190 3470
rect 19708 2060 19808 2070
rect 22130 2370 22230 2380
rect 19020 888 19120 1346
rect 19020 372 19120 830
rect 19020 -144 19120 314
rect 19020 -540 19120 -202
rect 21130 1970 21230 1980
rect 21130 1662 21230 1870
rect 21130 1146 21230 1604
rect 21130 630 21230 1088
rect 21130 114 21230 572
rect 21130 -402 21230 56
rect 21130 -540 21230 -460
rect 22130 1404 22230 2270
rect 23090 1970 23190 3090
rect 23550 2570 23650 2580
rect 23090 1860 23190 1870
rect 23390 2430 23490 2440
rect 22130 888 22230 1346
rect 22130 372 22230 830
rect 22130 -144 22230 314
rect 22130 -540 22230 -202
rect 23390 1662 23490 2330
rect 23390 1404 23490 1604
rect 23390 1146 23490 1346
rect 23390 888 23490 1088
rect 23390 630 23490 830
rect 23390 372 23490 572
rect 23390 114 23490 314
rect 23390 -144 23490 56
rect 23390 -402 23490 -202
rect 23390 -540 23490 -460
rect 23550 1570 23650 2470
rect 23620 1430 23650 1570
rect 23550 1320 23650 1430
rect 23620 1180 23650 1320
rect 23550 1060 23650 1180
rect 23620 920 23650 1060
rect 23550 800 23650 920
rect 23620 660 23650 800
rect 23550 550 23650 660
rect 23620 410 23650 550
rect 23550 290 23650 410
rect 23620 150 23650 290
rect 23550 30 23650 150
rect 23620 -110 23650 30
rect 23550 -230 23650 -110
rect 23620 -370 23650 -230
rect 23550 -540 23650 -370
<< via2 >>
rect 940 2470 1040 2570
rect 2738 2670 2838 2770
rect 4666 2470 4766 2570
rect 1140 2270 1240 2370
rect 3470 2270 3570 2370
rect 2470 1870 2570 1970
rect 6594 2270 6694 2370
rect 6800 2270 6900 2370
rect 13370 3720 13470 3820
rect 12378 2670 12478 2770
rect 10450 2470 10550 2570
rect 12800 2470 12900 2570
rect 8522 2270 8622 2370
rect 9690 2270 9790 2370
rect 5580 1870 5680 1970
rect 8690 1870 8790 1970
rect 16370 3730 16430 3830
rect 15720 3290 15820 3360
rect 15720 3260 15820 3290
rect 16460 3260 16560 3360
rect 16800 2670 16900 2770
rect 13920 2470 14020 2570
rect 13070 2270 13170 2370
rect 15910 2270 16010 2370
rect 14910 1870 15010 1970
rect 18288 2670 18388 2770
rect 18998 2670 19098 2770
rect 17578 2070 17678 2170
rect 19020 2270 19120 2370
rect 18020 1870 18120 1970
rect 20290 2670 20390 2770
rect 19708 2070 19808 2170
rect 22130 2270 22230 2370
rect 21130 1870 21230 1970
rect 23550 2470 23650 2570
rect 23090 1870 23190 1970
<< metal3 >>
rect 16360 3830 16440 3835
rect 13390 3825 16370 3830
rect 13360 3820 16370 3825
rect 13360 3720 13370 3820
rect 13470 3730 16370 3820
rect 16430 3730 16440 3830
rect 13470 3720 13480 3730
rect 16360 3725 16440 3730
rect 13360 3715 13480 3720
rect 15710 3360 15830 3365
rect 16450 3360 16570 3365
rect 15710 3260 15720 3360
rect 15820 3260 16460 3360
rect 16560 3260 16660 3360
rect 15710 3255 15830 3260
rect 16450 3255 16570 3260
rect 2728 2770 2848 2775
rect 12368 2770 12488 2775
rect 16790 2770 16910 2775
rect 18278 2770 18398 2775
rect 18988 2770 19108 2775
rect 20280 2770 20400 2775
rect 1280 2670 2738 2770
rect 2838 2670 12378 2770
rect 12478 2670 16800 2770
rect 16900 2670 18288 2770
rect 18388 2670 18998 2770
rect 19098 2670 20290 2770
rect 20390 2670 23520 2770
rect 2728 2665 2848 2670
rect 12368 2665 12488 2670
rect 16790 2665 16910 2670
rect 18278 2665 18398 2670
rect 18988 2665 19108 2670
rect 20280 2665 20400 2670
rect 930 2570 1050 2575
rect 4656 2570 4776 2575
rect 10440 2570 10560 2575
rect 12790 2570 12910 2575
rect 13910 2570 14030 2575
rect 23540 2570 23660 2575
rect 930 2470 940 2570
rect 1040 2470 4666 2570
rect 4766 2470 10450 2570
rect 10550 2470 12800 2570
rect 12900 2470 13920 2570
rect 14020 2470 23550 2570
rect 23650 2470 23660 2570
rect 930 2465 1050 2470
rect 4656 2465 4776 2470
rect 10440 2465 10560 2470
rect 12790 2465 12910 2470
rect 13910 2465 14030 2470
rect 23540 2465 23660 2470
rect 1130 2370 1250 2375
rect 3460 2370 3580 2375
rect 6584 2370 6704 2375
rect 6790 2370 6910 2375
rect 8512 2370 8632 2375
rect 9680 2370 9800 2375
rect 13060 2370 13180 2375
rect 15900 2370 16020 2375
rect 19010 2370 19130 2375
rect 22120 2370 22240 2375
rect 1130 2270 1140 2370
rect 1240 2270 3470 2370
rect 3570 2270 6594 2370
rect 6694 2270 6800 2370
rect 6900 2270 8522 2370
rect 8622 2270 9690 2370
rect 9790 2270 13070 2370
rect 13170 2270 15910 2370
rect 16010 2270 19020 2370
rect 19120 2270 22130 2370
rect 22230 2270 23520 2370
rect 1130 2265 1250 2270
rect 3460 2265 3580 2270
rect 6584 2265 6704 2270
rect 6790 2265 6910 2270
rect 8512 2265 8632 2270
rect 9680 2265 9800 2270
rect 13060 2265 13180 2270
rect 15900 2265 16020 2270
rect 19010 2265 19130 2270
rect 22120 2265 22240 2270
rect 17568 2170 17688 2175
rect 19698 2170 19818 2175
rect 1280 2070 17578 2170
rect 17678 2070 19708 2170
rect 19808 2070 23780 2170
rect 17568 2065 17688 2070
rect 19698 2065 19818 2070
rect 2460 1970 2580 1975
rect 5570 1970 5690 1975
rect 8680 1970 8800 1975
rect 14900 1970 15020 1975
rect 18010 1970 18130 1975
rect 21120 1970 21240 1975
rect 23080 1970 23200 1975
rect 1280 1870 2470 1970
rect 2570 1870 5580 1970
rect 5680 1870 8690 1970
rect 8790 1870 14910 1970
rect 15010 1870 18020 1970
rect 18120 1870 21130 1970
rect 21230 1870 23090 1970
rect 23190 1870 23520 1970
rect 2460 1865 2580 1870
rect 5570 1865 5690 1870
rect 8680 1865 8800 1870
rect 14900 1865 15020 1870
rect 18010 1865 18130 1870
rect 21120 1865 21240 1870
rect 23080 1865 23200 1870
use sky130_fd_pr__pfet_g5v0d10v5_8TN7ZV  XM1[1]
timestamp 1736799598
transform 0 1 6344 -1 0 3773
box -753 -1000 753 1000
use sky130_fd_pr__pfet_g5v0d10v5_8TN7ZV  XM1[2]
timestamp 1736799598
transform 0 -1 8272 1 0 3773
box -753 -1000 753 1000
use sky130_fd_pr__pfet_g5v0d10v5_8TN7ZV  XM2[1]
timestamp 1736799598
transform 0 1 4416 -1 0 3773
box -753 -1000 753 1000
use sky130_fd_pr__pfet_g5v0d10v5_8TN7ZV  XM2[2]
timestamp 1736799598
transform 0 1 10200 -1 0 3773
box -753 -1000 753 1000
use sky130_fd_pr__pfet_g5v0d10v5_8TN7ZV  XM3[1]
timestamp 1736799598
transform 0 1 12128 -1 0 3773
box -753 -1000 753 1000
use sky130_fd_pr__pfet_g5v0d10v5_8TN7ZV  XM3[2]
timestamp 1736799598
transform 0 1 2488 -1 0 3773
box -753 -1000 753 1000
use sky130_fd_pr__nfet_g5v0d10v5_T4FFC6  XM4[1]
timestamp 1736799799
transform 0 1 17528 -1 0 3757
box -687 -388 687 388
use sky130_fd_pr__nfet_g5v0d10v5_T4FFC6  XM4[2]
timestamp 1736799799
transform 0 1 19658 -1 0 3757
box -687 -388 687 388
use sky130_fd_pr__nfet_g5v0d10v5_T4FFC6  XM5[1]
timestamp 1736799799
transform 0 1 18238 -1 0 3757
box -687 -388 687 388
use sky130_fd_pr__nfet_g5v0d10v5_T4FFC6  XM5[2]
timestamp 1736799799
transform 0 1 18948 -1 0 3757
box -687 -388 687 388
use sky130_fd_pr__nfet_g5v0d10v5_Z9T923  XM6
timestamp 1736965693
transform 0 1 15028 1 0 3257
box -287 -1088 287 1088
use sky130_fd_pr__nfet_g5v0d10v5_NASXE7  XM7
timestamp 1736888431
transform -1 0 16528 0 -1 3878
box -158 -588 158 588
use sky130_fd_pr__pfet_g5v0d10v5_KH6JES  XM8
timestamp 1736888431
transform -1 0 14734 0 -1 4270
box -1124 -200 1124 200
use sky130_fd_pr__nfet_g5v0d10v5_8D664F  XM9
timestamp 1737184964
transform 0 1 12400 -1 0 601
box -1061 -1588 1061 1588
use sky130_fd_pr__nfet_g5v0d10v5_8D664F  XM10[1]
timestamp 1737184964
transform 0 1 3070 -1 0 601
box -1061 -1588 1061 1588
use sky130_fd_pr__nfet_g5v0d10v5_8D664F  XM10[2]
timestamp 1737184964
transform 0 1 6180 -1 0 601
box -1061 -1588 1061 1588
use sky130_fd_pr__nfet_g5v0d10v5_8D664F  XM10[3]
timestamp 1737184964
transform 0 1 9290 -1 0 601
box -1061 -1588 1061 1588
use sky130_fd_pr__nfet_g5v0d10v5_8D664F  XM10[4]
timestamp 1737184964
transform 0 1 15510 -1 0 601
box -1061 -1588 1061 1588
use sky130_fd_pr__nfet_g5v0d10v5_8D664F  XM10[5]
timestamp 1737184964
transform 0 1 18620 -1 0 601
box -1061 -1588 1061 1588
use sky130_fd_pr__nfet_g5v0d10v5_8D664F  XM10[6]
timestamp 1737184964
transform 0 1 21730 -1 0 601
box -1061 -1588 1061 1588
use sky130_fd_pr__pfet_g5v0d10v5_4DZKWV  XMDY1[1]
timestamp 1736799598
transform 0 -1 1360 1 0 3773
box -753 -200 753 200
use sky130_fd_pr__pfet_g5v0d10v5_9TWSB2  XMDY1[2]
timestamp 1736799799
transform 0 1 13256 -1 0 3773
box -753 -200 753 200
use sky130_fd_pr__nfet_g5v0d10v5_5XWZCB  XMDY2[1]
timestamp 1736799799
transform 0 1 17018 -1 0 3757
box -687 -188 687 188
use sky130_fd_pr__nfet_g5v0d10v5_5XWZCB  XMDY2[2]
timestamp 1736799799
transform 0 1 20168 -1 0 3757
box -687 -188 687 188
use sky130_fd_pr__nfet_g5v0d10v5_WC59T4  XMDY3[1]
timestamp 1737184964
transform 0 -1 23440 1 0 601
box -1061 -188 1061 188
use sky130_fd_pr__nfet_g5v0d10v5_WC59T4  XMDY3[2]
timestamp 1737184964
transform 0 1 1360 1 0 601
box -1061 -188 1061 188
use sky130_fd_pr__res_high_po_1p41_WUTXG4  XR1
timestamp 1737183131
transform 0 -1 21906 1 0 3708
box -708 -1446 708 1446
<< labels >>
flabel metal1 940 4880 1140 5080 0 FreeSans 256 180 0 0 vdda
port 0 nsew
flabel metal1 940 2530 1140 2730 0 FreeSans 256 180 0 0 vssa
port 2 nsew
flabel metal3 23680 2070 23780 2170 0 FreeSans 160 0 0 0 iptat
port 1 nsew
<< end >>
