magic
tech sky130A
magscale 1 2
timestamp 1736106420
<< nwell >>
rect -2540 6520 10420 7840
rect -2540 1810 8800 6520
<< mvpsubdiff >>
rect 8890 6310 10420 6430
rect 8890 1720 9010 6310
rect -2470 1600 9010 1720
rect -2470 840 -2350 1600
rect 10300 840 10420 6310
rect -2470 820 10420 840
rect -2470 740 2920 820
rect 3200 740 10420 820
rect -2470 720 10420 740
<< mvnsubdiff >>
rect -2470 7750 10350 7770
rect -2470 7670 -2070 7750
rect -1860 7670 10350 7750
rect -2470 7650 10350 7670
rect -2470 4870 -2350 7650
rect 8610 6710 8730 7650
rect 10230 6710 10350 7650
rect 8610 6590 10350 6710
rect 8610 4870 8730 6590
rect -2470 4750 8730 4870
rect -2470 2000 -2350 4750
rect 8610 2000 8730 4750
rect -2470 1880 8730 2000
<< mvpsubdiffcont >>
rect 2920 740 3200 820
<< mvnsubdiffcont >>
rect -2070 7670 -1860 7750
<< locali >>
rect -2450 7670 -2070 7750
rect -1860 7670 10330 7750
rect -2450 4850 -2370 7670
rect 8630 6690 8710 7670
rect 10250 6690 10330 7670
rect 8630 6610 10330 6690
rect 8630 4850 8710 6610
rect -2450 4770 8710 4850
rect -2450 1980 -2370 4770
rect 8630 1980 8710 4770
rect -2450 1900 8710 1980
rect 8910 6330 10400 6410
rect 8910 1700 8990 6330
rect -2450 1620 8990 1700
rect -2450 820 -2370 1620
rect 10320 820 10400 6330
rect -2450 740 2920 820
rect 3200 740 10400 820
<< viali >>
rect -2070 7670 -1860 7750
rect 2920 740 3200 820
<< metal1 >>
rect -2540 8020 10420 8050
rect -2540 8010 1476 8020
rect -2540 7850 -830 8010
rect -730 7850 98 8010
rect 198 7860 1476 8010
rect 1576 7860 2854 8020
rect 2954 7860 4232 8020
rect 4332 7860 5610 8020
rect 5710 7860 6988 8020
rect 7088 8010 10420 8020
rect 7088 7860 9490 8010
rect 198 7850 9490 7860
rect 9590 7850 10420 8010
rect -2540 7750 10420 7850
rect -2540 7670 -2070 7750
rect -1860 7670 10420 7750
rect -2540 7650 10420 7670
rect -2540 7640 -2330 7650
rect -840 7530 -830 7588
rect -730 7530 -720 7588
rect 88 7530 98 7588
rect 198 7530 208 7588
rect 1466 7530 1476 7588
rect 1576 7530 1586 7588
rect 2844 7530 2854 7588
rect 2954 7530 2964 7588
rect 4222 7530 4232 7588
rect 4332 7530 4342 7588
rect 5600 7530 5610 7588
rect 5710 7530 5720 7588
rect 6978 7530 6988 7588
rect 7088 7530 7098 7588
rect -990 7346 -980 7514
rect -910 7346 -900 7514
rect 7160 7346 7170 7514
rect 7240 7346 7250 7514
rect 9020 7402 9030 7530
rect 9090 7402 9100 7530
rect 9480 7516 9490 7574
rect 9590 7516 9600 7574
rect 9200 7358 9210 7416
rect 9310 7358 9320 7416
rect -840 7272 -830 7330
rect -730 7272 -720 7330
rect 538 7272 548 7330
rect 648 7272 658 7330
rect 1916 7272 1926 7330
rect 2026 7272 2036 7330
rect 3294 7272 3304 7330
rect 3404 7272 3414 7330
rect 4672 7272 4682 7330
rect 4782 7272 4792 7330
rect 6050 7272 6060 7330
rect 6160 7272 6170 7330
rect 6978 7272 6988 7330
rect 7088 7272 7098 7330
rect -990 7088 -980 7256
rect -910 7088 -900 7256
rect 7160 7088 7170 7256
rect 7240 7088 7250 7256
rect 9210 7080 9220 7250
rect 9280 7080 9290 7250
rect 9480 7224 9490 7282
rect 9590 7224 9600 7282
rect -840 7014 -830 7072
rect -730 7014 -720 7072
rect 88 7014 98 7072
rect 198 7014 208 7072
rect 1466 7014 1476 7072
rect 1576 7014 1586 7072
rect 2844 7014 2854 7072
rect 2954 7014 2964 7072
rect 4221 7014 4231 7072
rect 4331 7014 4341 7072
rect 5600 7014 5610 7072
rect 5710 7014 5720 7072
rect 6978 7014 6988 7072
rect 7088 7014 7098 7072
rect 9540 7066 9550 7124
rect 9650 7066 9660 7124
rect -990 6830 -980 6998
rect -910 6830 -900 6998
rect 7160 6830 7170 6998
rect 7240 6830 7250 6998
rect -840 6756 -830 6814
rect -730 6756 -720 6814
rect 538 6756 548 6814
rect 648 6756 658 6814
rect 1916 6756 1926 6814
rect 2026 6756 2036 6814
rect 3294 6756 3304 6814
rect 3404 6756 3414 6814
rect 4672 6756 4682 6814
rect 4782 6756 4792 6814
rect 6050 6756 6060 6814
rect 6160 6756 6170 6814
rect 6978 6756 6988 6814
rect 7088 6756 7098 6814
rect -990 6572 -980 6740
rect -910 6572 -900 6740
rect 7160 6572 7170 6740
rect 7240 6572 7250 6740
rect -840 6498 -830 6556
rect -730 6498 -720 6556
rect 88 6498 98 6556
rect 198 6498 208 6556
rect 1466 6498 1476 6556
rect 1576 6498 1586 6556
rect 2844 6498 2854 6556
rect 2954 6498 2964 6556
rect 4222 6498 4232 6556
rect 4332 6498 4342 6556
rect 5600 6498 5610 6556
rect 5710 6498 5720 6556
rect 6978 6498 6988 6556
rect 7088 6498 7098 6556
rect -990 6314 -980 6482
rect -910 6314 -900 6482
rect 7160 6314 7170 6482
rect 7240 6314 7250 6482
rect -840 6240 -830 6298
rect -730 6240 -720 6298
rect 538 6240 548 6298
rect 648 6240 658 6298
rect 1916 6240 1926 6298
rect 2026 6240 2036 6298
rect 3294 6240 3304 6298
rect 3404 6240 3414 6298
rect 4672 6240 4682 6298
rect 4782 6240 4792 6298
rect 6050 6240 6060 6298
rect 6160 6240 6170 6298
rect 6978 6240 6988 6298
rect 7088 6240 7098 6298
rect -990 6056 -980 6224
rect -910 6056 -900 6224
rect 7160 6056 7170 6224
rect 7240 6056 7250 6224
rect -840 5982 -830 6040
rect -730 5982 -720 6040
rect 88 5982 98 6040
rect 198 5982 208 6040
rect 1466 5982 1476 6040
rect 1576 5982 1586 6040
rect 2844 5982 2854 6040
rect 2954 5982 2964 6040
rect 4222 5982 4232 6040
rect 4332 5982 4342 6040
rect 5600 5982 5610 6040
rect 5710 5982 5720 6040
rect 6978 5982 6988 6040
rect 7088 5982 7098 6040
rect 9030 6010 9040 6160
rect 9100 6010 9110 6160
rect 9190 6128 9200 6186
rect 9320 6128 9330 6186
rect 9338 6134 9486 6180
rect 9440 6120 9486 6134
rect 9530 6128 9540 6186
rect 9660 6128 9670 6186
rect -990 5798 -980 5966
rect -910 5798 -900 5966
rect 7160 5798 7170 5966
rect 7240 5798 7250 5966
rect 9140 5900 10170 6000
rect 10270 5900 10280 6000
rect -840 5724 -830 5782
rect -730 5724 -720 5782
rect 538 5724 548 5782
rect 648 5724 658 5782
rect 1916 5724 1926 5782
rect 2026 5724 2036 5782
rect 3294 5724 3304 5782
rect 3404 5724 3414 5782
rect 4672 5724 4682 5782
rect 4782 5724 4792 5782
rect 6050 5724 6060 5782
rect 6160 5724 6170 5782
rect 6978 5724 6988 5782
rect 7088 5724 7098 5782
rect -990 5540 -980 5708
rect -910 5540 -900 5708
rect 7160 5540 7170 5708
rect 7240 5540 7250 5708
rect -840 5466 -830 5524
rect -730 5466 -720 5524
rect 88 5466 98 5524
rect 198 5466 208 5524
rect 1465 5466 1475 5524
rect 1575 5466 1585 5524
rect 2844 5466 2854 5524
rect 2954 5466 2964 5524
rect 4222 5465 4232 5523
rect 4332 5465 4342 5523
rect 5600 5466 5610 5524
rect 5710 5466 5720 5524
rect 6978 5466 6988 5524
rect 7088 5466 7098 5524
rect 9358 5330 9368 5430
rect 9426 5330 9436 5430
rect 9874 5330 9884 5430
rect 9942 5330 9952 5430
rect -1030 4634 -1020 4692
rect -920 4634 -910 4692
rect 2780 4640 2867 4686
rect 2821 4630 2867 4640
rect 3393 4640 3480 4686
rect 3393 4630 3439 4640
rect 7170 4634 7180 4692
rect 7280 4634 7290 4692
rect -1030 4376 -1020 4434
rect -920 4376 -910 4434
rect 7170 4376 7180 4434
rect 7280 4376 7290 4434
rect 2844 4226 2980 4326
rect 3080 4226 3090 4326
rect 220 4118 230 4176
rect 330 4118 340 4176
rect 2821 4080 2867 4180
rect 3393 4114 3439 4180
rect 5920 4118 5930 4176
rect 6030 4118 6040 4176
rect 3170 3968 3180 4068
rect 3280 3968 3416 4068
rect -1030 3860 -1020 3918
rect -920 3860 -910 3918
rect 7170 3860 7180 3918
rect 7280 3860 7290 3918
rect 2844 3710 3180 3810
rect 3280 3710 3290 3810
rect 1470 3602 1480 3660
rect 1580 3602 1590 3660
rect 2821 3598 2867 3664
rect 3393 3598 3439 3664
rect 4670 3602 4680 3660
rect 4780 3602 4790 3660
rect 2970 3452 2980 3552
rect 3080 3454 3416 3552
rect 3080 3452 3393 3454
rect -1030 3344 -1020 3402
rect -920 3344 -910 3402
rect 7170 3344 7180 3402
rect 7280 3344 7290 3402
rect 2844 3194 3180 3294
rect 3280 3194 3290 3294
rect 9100 3190 9110 3290
rect 9168 3190 9178 3290
rect 9616 3190 9626 3290
rect 9684 3190 9694 3290
rect 10132 3190 10142 3290
rect 10200 3190 10210 3290
rect 1470 3086 1480 3144
rect 1580 3086 1590 3144
rect 2821 3082 2867 3148
rect 3393 3082 3439 3148
rect 4670 3086 4680 3144
rect 4780 3086 4790 3144
rect 2970 2936 2980 3036
rect 3080 2938 3416 3036
rect 3080 2936 3393 2938
rect -1030 2828 -1020 2886
rect -920 2828 -910 2886
rect 7170 2828 7180 2886
rect 7280 2828 7290 2886
rect 2844 2678 2980 2778
rect 3080 2678 3090 2778
rect 220 2570 230 2628
rect 330 2570 340 2628
rect 2821 2566 2867 2632
rect 3393 2566 3439 2632
rect 5920 2570 5930 2628
rect 6030 2570 6040 2628
rect 3170 2420 3180 2520
rect 3280 2420 3416 2520
rect -1030 2312 -1020 2370
rect -920 2312 -910 2370
rect 7170 2312 7180 2370
rect 7280 2312 7290 2370
rect -1030 2054 -1020 2112
rect -920 2054 -910 2112
rect 2821 2106 2867 2153
rect 2780 2060 2867 2106
rect 3393 2106 3439 2143
rect 3393 2060 3489 2106
rect 7170 2054 7180 2112
rect 7280 2054 7290 2112
rect 9170 1920 9180 1990
rect 9360 1920 9370 1990
rect 9430 1920 9440 1990
rect 9620 1920 9630 1990
rect 9690 1920 9700 1990
rect 9880 1920 9890 1990
rect 9950 1920 9960 1990
rect 10140 1920 10150 1990
rect -1405 1446 -1395 1504
rect -1294 1446 -1284 1504
rect -95 1446 -85 1504
rect 16 1446 26 1504
rect 1815 1446 1825 1504
rect 1926 1446 1936 1504
rect 3725 1446 3735 1504
rect 3836 1446 3846 1504
rect 5635 1447 5645 1505
rect 5746 1447 5756 1505
rect 7545 1446 7555 1504
rect 7656 1446 7666 1504
rect -1740 1270 -1730 1420
rect -1670 1270 -1660 1420
rect 7920 1270 7930 1420
rect 7990 1270 8000 1420
rect -1405 1188 -1395 1246
rect -1294 1188 -1284 1246
rect 505 1188 515 1246
rect 615 1188 625 1246
rect 2415 1188 2425 1246
rect 2525 1188 2535 1246
rect 4324 1188 4334 1246
rect 4436 1188 4446 1246
rect 6234 1188 6244 1246
rect 6346 1188 6356 1246
rect 7545 1188 7555 1246
rect 7656 1188 7666 1246
rect -1740 1010 -1730 1160
rect -1670 1010 -1660 1160
rect 7920 1010 7930 1160
rect 7990 1010 8000 1160
rect -1405 930 -1395 988
rect -1294 930 -1284 988
rect -95 930 -85 988
rect 16 930 26 988
rect 1815 930 1825 988
rect 1926 930 1936 988
rect 3725 930 3735 988
rect 3836 930 3846 988
rect 5635 930 5645 988
rect 5746 930 5756 988
rect 7545 930 7555 988
rect 7656 930 7666 988
rect -2540 820 10420 840
rect -2540 740 2920 820
rect 3200 740 10420 820
rect -2540 640 10420 740
rect -2540 480 -1395 640
rect -1294 480 -85 640
rect 16 480 1825 640
rect 1926 480 3735 640
rect 3836 480 5645 640
rect 5746 480 7555 640
rect 7656 480 10170 640
rect 10270 480 10420 640
rect -2540 440 10420 480
<< via1 >>
rect -830 7850 -730 8010
rect 98 7850 198 8010
rect 1476 7860 1576 8020
rect 2854 7860 2954 8020
rect 4232 7860 4332 8020
rect 5610 7860 5710 8020
rect 6988 7860 7088 8020
rect 9490 7850 9590 8010
rect -830 7530 -730 7588
rect 98 7530 198 7588
rect 1476 7530 1576 7588
rect 2854 7530 2954 7588
rect 4232 7530 4332 7588
rect 5610 7530 5710 7588
rect 6988 7530 7088 7588
rect -980 7346 -910 7514
rect 7170 7346 7240 7514
rect 9030 7402 9090 7530
rect 9490 7516 9590 7574
rect 9210 7358 9310 7416
rect -830 7272 -730 7330
rect 548 7272 648 7330
rect 1926 7272 2026 7330
rect 3304 7272 3404 7330
rect 4682 7272 4782 7330
rect 6060 7272 6160 7330
rect 6988 7272 7088 7330
rect -980 7088 -910 7256
rect 7170 7088 7240 7256
rect 9220 7080 9280 7250
rect 9490 7224 9590 7282
rect -830 7014 -730 7072
rect 98 7014 198 7072
rect 1476 7014 1576 7072
rect 2854 7014 2954 7072
rect 4231 7014 4331 7072
rect 5610 7014 5710 7072
rect 6988 7014 7088 7072
rect 9550 7066 9650 7124
rect -980 6830 -910 6998
rect 7170 6830 7240 6998
rect -830 6756 -730 6814
rect 548 6756 648 6814
rect 1926 6756 2026 6814
rect 3304 6756 3404 6814
rect 4682 6756 4782 6814
rect 6060 6756 6160 6814
rect 6988 6756 7088 6814
rect -980 6572 -910 6740
rect 7170 6572 7240 6740
rect -830 6498 -730 6556
rect 98 6498 198 6556
rect 1476 6498 1576 6556
rect 2854 6498 2954 6556
rect 4232 6498 4332 6556
rect 5610 6498 5710 6556
rect 6988 6498 7088 6556
rect -980 6314 -910 6482
rect 7170 6314 7240 6482
rect -830 6240 -730 6298
rect 548 6240 648 6298
rect 1926 6240 2026 6298
rect 3304 6240 3404 6298
rect 4682 6240 4782 6298
rect 6060 6240 6160 6298
rect 6988 6240 7088 6298
rect -980 6056 -910 6224
rect 7170 6056 7240 6224
rect -830 5982 -730 6040
rect 98 5982 198 6040
rect 1476 5982 1576 6040
rect 2854 5982 2954 6040
rect 4232 5982 4332 6040
rect 5610 5982 5710 6040
rect 6988 5982 7088 6040
rect 9040 6010 9100 6160
rect 9200 6128 9320 6186
rect 9540 6128 9660 6186
rect -980 5798 -910 5966
rect 7170 5798 7240 5966
rect 10170 5900 10270 6000
rect -830 5724 -730 5782
rect 548 5724 648 5782
rect 1926 5724 2026 5782
rect 3304 5724 3404 5782
rect 4682 5724 4782 5782
rect 6060 5724 6160 5782
rect 6988 5724 7088 5782
rect -980 5540 -910 5708
rect 7170 5540 7240 5708
rect -830 5466 -730 5524
rect 98 5466 198 5524
rect 1475 5466 1575 5524
rect 2854 5466 2954 5524
rect 4232 5465 4332 5523
rect 5610 5466 5710 5524
rect 6988 5466 7088 5524
rect 9368 5330 9426 5430
rect 9884 5330 9942 5430
rect -1020 4634 -920 4692
rect 7180 4634 7280 4692
rect -1020 4376 -920 4434
rect 7180 4376 7280 4434
rect 2980 4226 3080 4326
rect 230 4118 330 4176
rect 5930 4118 6030 4176
rect 3180 3968 3280 4068
rect -1020 3860 -920 3918
rect 7180 3860 7280 3918
rect 3180 3710 3280 3810
rect 1480 3602 1580 3660
rect 4680 3602 4780 3660
rect 2980 3452 3080 3552
rect -1020 3344 -920 3402
rect 7180 3344 7280 3402
rect 3180 3194 3280 3294
rect 9110 3190 9168 3290
rect 9626 3190 9684 3290
rect 10142 3190 10200 3290
rect 1480 3086 1580 3144
rect 4680 3086 4780 3144
rect 2980 2936 3080 3036
rect -1020 2828 -920 2886
rect 7180 2828 7280 2886
rect 2980 2678 3080 2778
rect 230 2570 330 2628
rect 5930 2570 6030 2628
rect 3180 2420 3280 2520
rect -1020 2312 -920 2370
rect 7180 2312 7280 2370
rect -1020 2054 -920 2112
rect 7180 2054 7280 2112
rect 9180 1920 9360 1990
rect 9440 1920 9620 1990
rect 9700 1920 9880 1990
rect 9960 1920 10140 1990
rect -1395 1446 -1294 1504
rect -85 1446 16 1504
rect 1825 1446 1926 1504
rect 3735 1446 3836 1504
rect 5645 1447 5746 1505
rect 7555 1446 7656 1504
rect -1730 1270 -1670 1420
rect 7930 1270 7990 1420
rect -1395 1188 -1294 1246
rect 515 1188 615 1246
rect 2425 1188 2525 1246
rect 4334 1188 4436 1246
rect 6244 1188 6346 1246
rect 7555 1188 7656 1246
rect -1730 1010 -1670 1160
rect 7930 1010 7990 1160
rect -1395 930 -1294 988
rect -85 930 16 988
rect 1825 930 1926 988
rect 3735 930 3836 988
rect 5645 930 5746 988
rect 7555 930 7656 988
rect -1395 480 -1294 640
rect -85 480 16 640
rect 1825 480 1926 640
rect 3735 480 3836 640
rect 5645 480 5746 640
rect 7555 480 7656 640
rect 10170 480 10270 640
<< metal2 >>
rect 1476 8020 1576 8030
rect -830 8010 -730 8020
rect -994 7730 -894 7740
rect -994 7514 -894 7630
rect -994 7346 -980 7514
rect -910 7346 -894 7514
rect -994 7256 -894 7346
rect -994 7088 -980 7256
rect -910 7088 -894 7256
rect -994 6998 -894 7088
rect -994 6830 -980 6998
rect -910 6830 -894 6998
rect -994 6740 -894 6830
rect -994 6572 -980 6740
rect -910 6572 -894 6740
rect -994 6482 -894 6572
rect -994 6314 -980 6482
rect -910 6314 -894 6482
rect -994 6224 -894 6314
rect -994 6056 -980 6224
rect -910 6056 -894 6224
rect -994 5966 -894 6056
rect -994 5798 -980 5966
rect -910 5798 -894 5966
rect -994 5708 -894 5798
rect -994 5540 -980 5708
rect -910 5540 -894 5708
rect -994 5430 -894 5540
rect -830 7588 -730 7850
rect -830 7330 -730 7530
rect -830 7072 -730 7272
rect -830 6814 -730 7014
rect -830 6556 -730 6756
rect -830 6298 -730 6498
rect -830 6040 -730 6240
rect -830 5782 -730 5982
rect -830 5524 -730 5724
rect -830 5430 -730 5466
rect 98 8010 198 8020
rect 98 7588 198 7850
rect 98 7072 198 7530
rect 98 6556 198 7014
rect 98 6040 198 6498
rect 98 5524 198 5982
rect 98 5430 198 5466
rect 548 7330 648 7624
rect 548 6814 648 7272
rect 548 6298 648 6756
rect 548 5782 648 6240
rect -1020 5230 -920 5240
rect -1020 4692 -920 5130
rect 548 5230 648 5724
rect 1476 7588 1576 7860
rect 2854 8020 2954 8030
rect 1476 7072 1576 7530
rect 1476 6556 1576 7014
rect 1476 6040 1576 6498
rect 1476 5534 1576 5982
rect 1475 5524 1576 5534
rect 1575 5466 1576 5524
rect 1475 5456 1576 5466
rect 1476 5430 1576 5456
rect 1926 7330 2026 7624
rect 1926 6814 2026 7272
rect 1926 6298 2026 6756
rect 1926 5782 2026 6240
rect 1926 5440 2026 5724
rect 2854 7588 2954 7860
rect 4232 8020 4332 8030
rect 2854 7072 2954 7530
rect 2854 6556 2954 7014
rect 2854 6040 2954 6498
rect 2854 5524 2954 5982
rect 1926 5430 2027 5440
rect 2854 5430 2954 5466
rect 3304 7730 3404 7740
rect 3304 7330 3404 7630
rect 3304 6814 3404 7272
rect 4232 7588 4332 7860
rect 5610 8020 5710 8030
rect 4232 7082 4332 7530
rect 4231 7072 4332 7082
rect 4331 7014 4332 7072
rect 4231 7004 4332 7014
rect 3304 6298 3404 6756
rect 3304 5782 3404 6240
rect 3304 5430 3404 5724
rect 4232 6556 4332 7004
rect 4232 6040 4332 6498
rect 4232 5523 4332 5982
rect 4232 5430 4332 5465
rect 4682 7330 4782 7624
rect 4682 6814 4782 7272
rect 4682 6298 4782 6756
rect 4682 5782 4782 6240
rect 4682 5430 4782 5724
rect 5610 7588 5710 7860
rect 6988 8020 7088 8030
rect 5610 7072 5710 7530
rect 5610 6556 5710 7014
rect 5610 6040 5710 6498
rect 5610 5524 5710 5982
rect 5610 5430 5710 5466
rect 6060 7330 6160 7624
rect 6060 6814 6160 7272
rect 6060 6298 6160 6756
rect 6060 5782 6160 6240
rect 1926 5320 2027 5330
rect 4682 5320 4782 5330
rect 548 5120 648 5130
rect 6060 5230 6160 5724
rect 6988 7588 7088 7860
rect 9490 8010 9590 8020
rect 6988 7330 7088 7530
rect 6988 7072 7088 7272
rect 6988 6814 7088 7014
rect 6988 6556 7088 6756
rect 6988 6298 7088 6498
rect 6988 6040 7088 6240
rect 6988 5782 7088 5982
rect 6988 5524 7088 5724
rect 6988 5430 7088 5466
rect 7152 7730 7252 7740
rect 7152 7514 7252 7630
rect 9490 7574 9590 7850
rect 7152 7346 7170 7514
rect 7240 7346 7252 7514
rect 7152 7256 7252 7346
rect 7152 7088 7170 7256
rect 7240 7088 7252 7256
rect 7152 6998 7252 7088
rect 7152 6830 7170 6998
rect 7240 6830 7252 6998
rect 7152 6740 7252 6830
rect 7152 6572 7170 6740
rect 7240 6572 7252 6740
rect 7152 6482 7252 6572
rect 7152 6314 7170 6482
rect 7240 6314 7252 6482
rect 7152 6224 7252 6314
rect 7152 6056 7170 6224
rect 7240 6056 7252 6224
rect 7152 5966 7252 6056
rect 7152 5798 7170 5966
rect 7240 5798 7252 5966
rect 7152 5708 7252 5798
rect 7152 5540 7170 5708
rect 7240 5540 7252 5708
rect 7152 5430 7252 5540
rect 9010 7530 9110 7540
rect 9010 7402 9030 7530
rect 9090 7402 9110 7530
rect 9010 6160 9110 7402
rect 9210 7416 9310 7426
rect 9210 7250 9310 7358
rect 9210 7080 9220 7250
rect 9280 7080 9310 7250
rect 9490 7282 9590 7516
rect 9490 7214 9590 7224
rect 9210 6196 9310 7080
rect 9550 7124 9650 7134
rect 9550 6310 9650 7066
rect 9550 6196 9650 6210
rect 9010 6010 9040 6160
rect 9100 6010 9110 6160
rect 9200 6186 9320 6196
rect 9200 6118 9320 6128
rect 9540 6186 9660 6196
rect 9540 6118 9660 6128
rect 9010 5430 9110 6010
rect 10170 6000 10270 6010
rect 9010 5320 9110 5330
rect 9368 5430 9426 5440
rect 9368 5320 9426 5330
rect 9884 5430 9942 5440
rect 9884 5320 9942 5330
rect 6060 5120 6160 5130
rect 7180 5230 7280 5240
rect 3180 5030 3280 5040
rect 2980 4830 3080 4840
rect -1020 4434 -920 4634
rect -1020 3918 -920 4376
rect -1020 3402 -920 3860
rect -1020 2886 -920 3344
rect -1020 2370 -920 2828
rect -1020 2112 -920 2312
rect -1020 2020 -920 2054
rect 230 4176 330 4690
rect 230 2628 330 4118
rect -1750 1820 -1650 1830
rect -1750 1420 -1650 1720
rect 230 1820 330 2570
rect 1480 3660 1580 4700
rect 1480 3144 1580 3602
rect 230 1710 330 1720
rect 515 2020 615 2030
rect -1750 1270 -1730 1420
rect -1670 1270 -1650 1420
rect -1750 1160 -1650 1270
rect -1750 1010 -1730 1160
rect -1670 1010 -1650 1160
rect -1750 930 -1650 1010
rect -1395 1504 -1294 1514
rect -1395 1436 -1294 1446
rect -85 1504 16 1514
rect -85 1436 16 1446
rect -1395 1256 -1295 1436
rect -1395 1246 -1294 1256
rect -1395 1178 -1294 1188
rect -1395 998 -1295 1178
rect -85 998 15 1436
rect 515 1246 615 1920
rect 1480 2020 1580 3086
rect 2980 4326 3080 4730
rect 2980 3552 3080 4226
rect 2980 3036 3080 3452
rect 2980 2778 3080 2936
rect 2980 2020 3080 2678
rect 3180 4068 3280 4930
rect 3180 3810 3280 3968
rect 3180 3294 3280 3710
rect 3180 2520 3280 3194
rect 3180 2020 3280 2420
rect 4680 3660 4780 4700
rect 4680 3144 4780 3602
rect 1480 1910 1580 1920
rect 2425 1820 2525 1830
rect -1395 988 -1294 998
rect -1395 920 -1294 930
rect -85 988 16 998
rect -1395 650 -1295 920
rect -1395 640 -1294 650
rect -1395 470 -1294 480
rect -85 640 16 930
rect 515 920 615 1188
rect 1825 1504 1926 1514
rect 1825 1436 1926 1446
rect 1825 998 1925 1436
rect 2425 1246 2525 1720
rect 4335 1820 4435 1830
rect 1825 988 1926 998
rect -85 470 16 480
rect 1825 640 1926 930
rect 2425 920 2525 1188
rect 3735 1504 3836 1514
rect 3735 1436 3836 1446
rect 3735 998 3835 1436
rect 4335 1256 4435 1720
rect 4680 1820 4780 3086
rect 5930 4176 6030 4700
rect 5930 2628 6030 4118
rect 5930 2020 6030 2570
rect 7180 4692 7280 5130
rect 7180 4434 7280 4634
rect 7180 3918 7280 4376
rect 7180 3402 7280 3860
rect 7180 2886 7280 3344
rect 10170 3300 10270 5900
rect 9110 3290 9168 3300
rect 9110 3180 9168 3190
rect 9626 3290 9684 3300
rect 9626 3180 9684 3190
rect 10142 3290 10270 3300
rect 10200 3190 10270 3290
rect 10142 3180 10270 3190
rect 7180 2370 7280 2828
rect 7180 2112 7280 2312
rect 7180 2044 7280 2054
rect 5930 1910 6030 1920
rect 6245 2020 6345 2030
rect 4680 1710 4780 1720
rect 5645 1505 5746 1515
rect 5645 1437 5746 1447
rect 4334 1246 4436 1256
rect 4334 1178 4436 1188
rect 3735 988 3836 998
rect 1825 470 1926 480
rect 3735 640 3836 930
rect 4335 920 4435 1178
rect 5645 998 5745 1437
rect 6245 1256 6345 1920
rect 9180 1990 9360 2000
rect 9180 1910 9360 1920
rect 9440 1990 9620 2000
rect 9440 1910 9620 1920
rect 9700 1990 9880 2000
rect 9700 1910 9880 1920
rect 9960 1990 10140 2000
rect 9960 1910 10140 1920
rect 7910 1820 8010 1830
rect 7555 1504 7656 1514
rect 7555 1436 7656 1446
rect 7555 1256 7655 1436
rect 7910 1420 8010 1720
rect 7910 1270 7930 1420
rect 7990 1270 8010 1420
rect 6244 1246 6346 1256
rect 6244 1178 6346 1188
rect 7555 1246 7656 1256
rect 7555 1178 7656 1188
rect 5645 988 5746 998
rect 3735 470 3836 480
rect 5645 640 5746 930
rect 6245 920 6345 1178
rect 7555 998 7655 1178
rect 7910 1160 8010 1270
rect 7910 1010 7930 1160
rect 7990 1010 8010 1160
rect 7555 988 7656 998
rect 7910 930 8010 1010
rect 5645 470 5746 480
rect 7555 640 7656 930
rect 7555 470 7656 480
rect 10170 640 10270 3180
rect 10170 470 10270 480
<< via2 >>
rect -994 7630 -894 7730
rect -1020 5130 -920 5230
rect 3304 7630 3404 7730
rect 1926 5330 2027 5430
rect 4682 5330 4782 5430
rect 548 5130 648 5230
rect 7152 7630 7252 7730
rect 9550 6210 9650 6310
rect 9010 5330 9110 5430
rect 9368 5330 9426 5430
rect 9884 5330 9942 5430
rect 6060 5130 6160 5230
rect 7180 5130 7280 5230
rect 3180 4930 3280 5030
rect 2980 4730 3080 4830
rect -1750 1720 -1650 1820
rect 230 1720 330 1820
rect 515 1920 615 2020
rect 1480 1920 1580 2020
rect 2425 1720 2525 1820
rect 4335 1720 4435 1820
rect 9110 3190 9168 3290
rect 9626 3190 9684 3290
rect 10142 3190 10200 3290
rect 5930 1920 6030 2020
rect 6245 1920 6345 2020
rect 4680 1720 4780 1820
rect 9180 1920 9360 1990
rect 9440 1920 9620 1990
rect 9700 1920 9880 1990
rect 9960 1920 10140 1990
rect 7910 1720 8010 1820
<< metal3 >>
rect -1004 7730 -884 7735
rect 3294 7730 3414 7735
rect 7142 7730 7262 7735
rect -2540 7630 -994 7730
rect -894 7630 3304 7730
rect 3404 7630 7152 7730
rect 7252 7630 7262 7730
rect -1004 7625 -884 7630
rect 3294 7625 3414 7630
rect 7142 7625 7262 7630
rect 9540 6310 9660 6315
rect 9540 6210 9550 6310
rect 9650 6210 10420 6310
rect 9540 6205 9660 6210
rect 1916 5430 2037 5435
rect 4672 5430 4792 5435
rect 9000 5430 9120 5435
rect 9358 5430 9436 5435
rect 9874 5430 9952 5435
rect -860 5330 1926 5430
rect 2027 5330 4682 5430
rect 4782 5330 9010 5430
rect 9110 5330 9368 5430
rect 9426 5330 9884 5430
rect 9942 5330 10210 5430
rect 1916 5325 2037 5330
rect 4672 5325 4792 5330
rect 9000 5325 9120 5330
rect 9358 5325 9436 5330
rect 9874 5325 9952 5330
rect -1030 5230 -910 5235
rect 538 5230 658 5235
rect 6050 5230 6170 5235
rect 7170 5230 7290 5235
rect -2400 5130 -1020 5230
rect -920 5130 548 5230
rect 648 5130 6060 5230
rect 6160 5130 7180 5230
rect 7280 5130 8600 5230
rect -1030 5125 -910 5130
rect 538 5125 658 5130
rect 6050 5125 6170 5130
rect 7170 5125 7290 5130
rect 3170 5030 3290 5035
rect -2540 4930 3180 5030
rect 3280 4930 8600 5030
rect 3170 4925 3290 4930
rect 2970 4830 3090 4835
rect -2540 4730 2980 4830
rect 3080 4730 8600 4830
rect 2970 4725 3090 4730
rect 9100 3290 9178 3295
rect 9616 3290 9694 3295
rect 10132 3290 10210 3295
rect 9100 3190 9110 3290
rect 9168 3190 9626 3290
rect 9684 3190 10142 3290
rect 10200 3190 10240 3290
rect 9100 3185 9178 3190
rect 9616 3185 9694 3190
rect 10132 3185 10210 3190
rect 505 2020 625 2025
rect 1470 2020 1590 2025
rect 5920 2020 6040 2025
rect 6235 2020 6355 2025
rect -2320 1920 515 2020
rect 615 1920 1480 2020
rect 1580 1920 5930 2020
rect 6030 1920 6245 2020
rect 6345 1990 10200 2020
rect 6345 1920 9180 1990
rect 9360 1920 9440 1990
rect 9620 1920 9700 1990
rect 9880 1920 9960 1990
rect 10140 1920 10200 1990
rect 505 1915 625 1920
rect 1470 1915 1590 1920
rect 5920 1915 6040 1920
rect 6235 1915 6355 1920
rect 9170 1915 9370 1920
rect 9430 1915 9630 1920
rect 9690 1915 9890 1920
rect 9950 1915 10150 1920
rect -1760 1820 -1640 1825
rect 220 1820 340 1825
rect 2415 1820 2535 1825
rect 4325 1820 4445 1825
rect 4670 1820 4790 1825
rect 7900 1820 8020 1825
rect -2320 1720 -1750 1820
rect -1650 1720 230 1820
rect 330 1720 2425 1820
rect 2525 1720 4335 1820
rect 4435 1720 4680 1820
rect 4780 1720 7910 1820
rect 8010 1720 8580 1820
rect -1760 1715 -1640 1720
rect 220 1715 340 1720
rect 2415 1715 2535 1720
rect 4325 1715 4445 1720
rect 4670 1715 4790 1720
rect 7900 1715 8020 1720
use sky130_fd_pr__pfet_g5v0d10v5_WRFAJJ  XM1[1]
timestamp 1736061100
transform 0 -1 373 -1 0 6527
box -1127 -725 1127 725
use sky130_fd_pr__pfet_g5v0d10v5_WRFAJJ  XM1[2]
timestamp 1736061100
transform 0 1 5885 -1 0 6527
box -1127 -725 1127 725
use sky130_fd_pr__pfet_g5v0d10v5_WRFAJJ  XM2
timestamp 1736061100
transform 0 1 3129 -1 0 6527
box -1127 -725 1127 725
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM3[1]
timestamp 1735905531
transform 0 1 280 -1 0 4147
box -353 -2600 353 2600
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM3[2]
timestamp 1735905531
transform 0 1 5980 -1 0 3631
box -353 -2600 353 2600
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM3[3]
timestamp 1735905531
transform 0 1 5980 -1 0 3115
box -353 -2600 353 2600
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM3[4]
timestamp 1735905531
transform 0 1 280 -1 0 2599
box -353 -2600 353 2600
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM4[1]
timestamp 1735905531
transform 0 1 5980 1 0 4147
box -353 -2600 353 2600
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM4[2]
timestamp 1735905531
transform 0 -1 280 -1 0 3631
box -353 -2600 353 2600
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM4[3]
timestamp 1735905531
transform 0 -1 280 -1 0 3115
box -353 -2600 353 2600
use sky130_fd_pr__pfet_g5v0d10v5_JS2SSJ  XM4[4]
timestamp 1735905531
transform 0 -1 5980 -1 0 2599
box -353 -2600 353 2600
use sky130_fd_pr__nfet_g5v0d10v5_697GFE  XM5[1]
timestamp 1735905635
transform 0 1 265 -1 0 1217
box -287 -988 287 988
use sky130_fd_pr__nfet_g5v0d10v5_697GFE  XM5[2]
timestamp 1735905635
transform 0 -1 5995 -1 0 1217
box -287 -988 287 988
use sky130_fd_pr__nfet_g5v0d10v5_697GFE  XM6[1]
timestamp 1735905635
transform 0 1 2175 -1 0 1217
box -287 -988 287 988
use sky130_fd_pr__nfet_g5v0d10v5_697GFE  XM6[2]
timestamp 1735905635
transform 0 1 4085 1 0 1217
box -287 -988 287 988
use sky130_fd_pr__pfet_g5v0d10v5_KSGYUE  XM7
timestamp 1736080880
transform 0 1 9584 -1 0 7174
box -174 -364 174 402
use sky130_fd_pr__nfet_g5v0d10v5_SMV9TY  XM8
timestamp 1736080880
transform 0 -1 9587 -1 0 6078
box -108 -157 108 157
use sky130_fd_pr__nfet_g5v0d10v5_233RRQ  XM9
timestamp 1735905635
transform 1 0 9655 0 1 3768
box -545 -1838 545 1838
use sky130_fd_pr__pfet_g5v0d10v5_WRFAJJ  XM10[1]
timestamp 1736061100
transform 0 1 1751 -1 0 6527
box -1127 -725 1127 725
use sky130_fd_pr__pfet_g5v0d10v5_WRFAJJ  XM10[2]
timestamp 1736061100
transform 0 1 4507 -1 0 6527
box -1127 -725 1127 725
use sky130_fd_pr__pfet_g5v0d10v5_PE3VUG  XM11
timestamp 1736080880
transform 0 -1 9392 -1 0 7466
box -174 -402 174 364
use sky130_fd_pr__nfet_g5v0d10v5_SMV9TY  XM12
timestamp 1736080880
transform 0 -1 9207 1 0 6078
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_EWLYZD  XMDY1[1]
timestamp 1735905388
transform 0 1 -630 -1 0 6527
box -1127 -350 1127 350
use sky130_fd_pr__pfet_g5v0d10v5_EWLYZD  XMDY1[2]
timestamp 1735905388
transform 0 1 6888 -1 0 6527
box -1127 -350 1127 350
use sky130_fd_pr__pfet_g5v0d10v5_JSWDFN  XMDY2[1]
timestamp 1735905531
transform 0 1 280 -1 0 4534
box -224 -2600 224 2600
use sky130_fd_pr__pfet_g5v0d10v5_JSWDFN  XMDY2[2]
timestamp 1735905531
transform 0 1 5980 1 0 4534
box -224 -2600 224 2600
use sky130_fd_pr__pfet_g5v0d10v5_JSWDFN  XMDY2[3]
timestamp 1735905531
transform 0 -1 280 -1 0 2212
box -224 -2600 224 2600
use sky130_fd_pr__pfet_g5v0d10v5_JSWDFN  XMDY2[4]
timestamp 1735905531
transform 0 1 5980 -1 0 2212
box -224 -2600 224 2600
use sky130_fd_pr__nfet_g5v0d10v5_HEHGAL  XMDY3[1]
timestamp 1735905635
transform 0 1 -1195 -1 0 1217
box -287 -538 287 538
use sky130_fd_pr__nfet_g5v0d10v5_HEHGAL  XMDY3[2]
timestamp 1735905635
transform 0 1 7455 -1 0 1217
box -287 -538 287 538
<< labels >>
flabel metal3 10320 6210 10420 6310 0 FreeSans 160 0 0 0 outp
port 11 nsew
flabel metal3 -2540 4930 -2440 5030 0 FreeSans 160 0 0 0 inp
port 3 nsew
flabel metal3 -2540 4730 -2440 4830 0 FreeSans 160 0 0 0 inn
port 2 nsew
flabel metal1 -2540 440 -2340 640 0 FreeSans 256 180 0 0 vssa
port 5 nsew
flabel metal1 -2540 7850 -2340 8050 0 FreeSans 256 180 0 0 vdda
port 0 nsew
flabel metal3 -2540 7630 -2440 7730 0 FreeSans 160 0 0 0 ibias
port 1 nsew
<< end >>
