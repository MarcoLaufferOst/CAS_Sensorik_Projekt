* NGSPICE file created from r2r_dac_parax.ext - technology: sky130A

.subckt r2r_dac_parax V_out D1 D2 D5 D7 D4 V_REF D6 D3 D0 V_COM
X0 V_REF.t43 D1.t0 R2R_20k_0.B1.t1 V_REF.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X1 R2R_20k_0.B1.t6 a_372_n2638# V_COM.t69 sky130_fd_pr__res_xhigh_po_0p69 l=7
X2 R2R_20k_0.B0.t6 D0.t0 V_REF.t15 V_REF.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X3 V_REF.t9 D5.t0 R2R_20k_0.B5.t5 V_REF.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X4 R2R_20k_0.B1.t0 D1.t1 V_COM.t64 V_COM.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X5 R2R_20k_0.B7.t3 D7.t0 V_COM.t40 V_COM.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X6 R2R_20k_0.B6.t5 a_3882_n2638# V_COM.t38 sky130_fd_pr__res_xhigh_po_0p69 l=7
X7 R2R_20k_0.B4.t6 D4.t0 V_REF.t11 V_REF.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X8 V_REF.t37 D4.t1 R2R_20k_0.B4.t5 V_REF.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X9 a_1542_n838# a_1776_n2638# V_COM.t33 sky130_fd_pr__res_xhigh_po_0p69 l=7
X10 R2R_20k_0.B2.t5 D2.t0 V_REF.t25 V_REF.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X11 R2R_20k_0.B2.t2 D2.t1 V_COM.t75 V_COM.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X12 a_138_n838# a_n564_n838# V_COM.t47 sky130_fd_pr__res_xhigh_po_0p69 l=7
X13 R2R_20k_0.B6.t4 D6.t0 V_REF.t27 V_REF.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X14 R2R_20k_0.B2.t1 D2.t2 V_COM.t20 V_COM.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X15 R2R_20k_0.B7.t2 D7.t1 V_COM.t52 V_COM.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X16 a_2946_n838# a_3180_n2638# V_COM.t50 sky130_fd_pr__res_xhigh_po_0p69 l=7
X17 R2R_20k_0.B6.t2 D6.t1 V_REF.t17 V_REF.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X18 a_1542_n838# a_840_n838# V_COM.t46 sky130_fd_pr__res_xhigh_po_0p69 l=7
X19 R2R_20k_0.B5.t4 D5.t1 V_REF.t21 V_REF.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X20 V_REF.t47 D7.t2 R2R_20k_0.B7.t6 V_REF.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X21 a_3648_n838# a_2946_n838# V_COM.t66 sky130_fd_pr__res_xhigh_po_0p69 l=7
X22 R2R_20k_0.B0.t5 D0.t1 V_REF.t23 V_REF.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X23 R2R_20k_0.B3.t3 D3.t0 V_COM.t24 V_COM.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X24 a_840_n838# a_1074_n2638# V_COM.t73 sky130_fd_pr__res_xhigh_po_0p69 l=7
X25 V_COM.t71 V_COM.t72 V_COM.t70 sky130_fd_pr__res_xhigh_po_0p69 l=7
X26 R2R_20k_0.B3.t6 D3.t1 V_REF.t3 V_REF.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X27 V_REF.t33 D6.t2 R2R_20k_0.B6.t6 V_REF.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X28 V_COM.t77 V_COM.t78 V_COM.t76 sky130_fd_pr__res_xhigh_po_0p69 l=7
X29 V_COM.t68 a_n798_n2638# V_COM.t67 sky130_fd_pr__res_xhigh_po_0p69 l=7
X30 R2R_20k_0.B5.t6 a_3180_n2638# V_COM.t79 sky130_fd_pr__res_xhigh_po_0p69 l=7
X31 R2R_20k_0.B1.t2 D1.t2 V_REF.t41 V_REF.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X32 R2R_20k_0.B3.t2 D3.t2 V_COM.t7 V_COM.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X33 R2R_20k_0.B4.t3 D4.t2 V_COM.t18 V_COM.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X34 R2R_20k_0.B1.t3 D1.t3 V_REF.t39 V_REF.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X35 R2R_20k_0.B0.t3 D0.t2 V_COM.t12 V_COM.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X36 V_COM.t32 D5.t2 R2R_20k_0.B5.t2 V_COM.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X37 V_COM.t56 D4.t3 R2R_20k_0.B4.t2 V_COM.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X38 R2R_20k_0.B7.t5 D7.t3 V_REF.t29 V_REF.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X39 R2R_20k_0.B1.t4 D1.t4 V_COM.t62 V_COM.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X40 R2R_20k_0.B6.t3 D6.t3 V_COM.t27 V_COM.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X41 a_n564_n838# a_n798_n2638# V_COM.t58 sky130_fd_pr__res_xhigh_po_0p69 l=7
X42 V_REF.t7 D0.t3 R2R_20k_0.B0.t4 V_REF.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X43 R2R_20k_0.B5.t3 D5.t3 V_REF.t19 V_REF.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X44 V_COM.t29 D3.t3 R2R_20k_0.B3.t1 V_COM.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X45 R2R_20k_0.B5.t1 D5.t4 V_COM.t49 V_COM.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X46 R2R_20k_0.B2.t6 a_1074_n2638# V_COM.t65 sky130_fd_pr__res_xhigh_po_0p69 l=7
X47 V_out.t1 a_4584_n2638# V_COM.t57 sky130_fd_pr__res_xhigh_po_0p69 l=7
X48 V_REF.t13 D2.t3 R2R_20k_0.B2.t4 V_REF.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X49 R2R_20k_0.B0.t2 D0.t4 V_COM.t10 V_COM.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X50 R2R_20k_0.B4.t1 D4.t4 V_COM.t16 V_COM.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=2.03 pd=14.58 as=1.015 ps=7.29 w=7 l=0.5
X51 a_840_n838# a_138_n838# V_COM.t43 sky130_fd_pr__res_xhigh_po_0p69 l=7
X52 a_2946_n838# a_2244_n838# V_COM.t41 sky130_fd_pr__res_xhigh_po_0p69 l=7
X53 V_COM.t54 D0.t5 R2R_20k_0.B0.t1 V_COM.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X54 R2R_20k_0.B5.t0 D5.t5 V_COM.t45 V_COM.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X55 V_out.t0 a_3648_n838# V_COM.t5 sky130_fd_pr__res_xhigh_po_0p69 l=7
X56 V_COM.t60 D1.t5 R2R_20k_0.B1.t5 V_COM.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X57 a_2244_n838# a_2478_n2638# V_COM.t37 sky130_fd_pr__res_xhigh_po_0p69 l=7
X58 R2R_20k_0.B4.t0 a_2478_n2638# V_COM.t4 sky130_fd_pr__res_xhigh_po_0p69 l=7
X59 R2R_20k_0.B2.t3 D2.t4 V_REF.t5 V_REF.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=4.64 pd=32.58 as=2.32 ps=16.29 w=16 l=0.5
X60 a_138_n838# a_372_n2638# V_COM.t30 sky130_fd_pr__res_xhigh_po_0p69 l=7
X61 R2R_20k_0.B7.t4 D7.t4 V_REF.t31 V_REF.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X62 R2R_20k_0.B7.t0 a_4584_n2638# V_COM.t25 sky130_fd_pr__res_xhigh_po_0p69 l=7
X63 R2R_20k_0.B4.t4 D4.t5 V_REF.t45 V_REF.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X64 a_n564_n838# a_n330_n2638# V_COM.t36 sky130_fd_pr__res_xhigh_po_0p69 l=7
X65 a_2244_n838# a_1542_n838# V_COM.t3 sky130_fd_pr__res_xhigh_po_0p69 l=7
X66 V_REF.t1 D3.t4 R2R_20k_0.B3.t5 V_REF.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=2.32 ps=16.29 w=16 l=0.5
X67 R2R_20k_0.B6.t1 D6.t4 V_COM.t22 V_COM.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=2.03 ps=14.58 w=7 l=0.5
X68 R2R_20k_0.B3.t4 D3.t5 V_REF.t35 V_REF.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32 pd=16.29 as=4.64 ps=32.58 w=16 l=0.5
X69 R2R_20k_0.B0.t0 a_n330_n2638# V_COM.t2 sky130_fd_pr__res_xhigh_po_0p69 l=7
X70 a_3648_n838# a_3882_n2638# V_COM.t8 sky130_fd_pr__res_xhigh_po_0p69 l=7
X71 V_COM.t14 D2.t5 R2R_20k_0.B2.t0 V_COM.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X72 V_COM.t1 D6.t5 R2R_20k_0.B6.t0 V_COM.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X73 V_COM.t35 D7.t5 R2R_20k_0.B7.t1 V_COM.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=1.015 pd=7.29 as=1.015 ps=7.29 w=7 l=0.5
X74 R2R_20k_0.B3.t0 a_1776_n2638# V_COM.t42 sky130_fd_pr__res_xhigh_po_0p69 l=7
R0 D1.n5 D1.t3 963.587
R1 D1.n0 D1.t0 963.587
R2 D1.n1 D1.t2 963.587
R3 D1.n2 D1.t1 515.91
R4 D1.n3 D1.t5 515.91
R5 D1.n4 D1.t4 515.91
R6 D1.n4 D1.n3 59.4829
R7 D1.n3 D1.n2 59.4829
R8 D1.n3 D1.n0 9.54099
R9 D1.n5 D1.n4 9.54099
R10 D1.n2 D1.n1 9.54099
R11 D1 D1.n6 7.56993
R12 D1 D1.n0 0.063
R13 D1.n6 D1.n5 0.0604957
R14 D1.n6 D1.n0 0.0402155
R15 D1.n1 D1 0.03675
R16 R2R_20k_0.B1.n5 R2R_20k_0.B1.t6 21.7027
R17 R2R_20k_0.B1.n3 R2R_20k_0.B1.t3 20.8848
R18 R2R_20k_0.B1.n2 R2R_20k_0.B1.n0 19.1576
R19 R2R_20k_0.B1.n3 R2R_20k_0.B1.t4 12.3059
R20 R2R_20k_0.B1.n2 R2R_20k_0.B1.n1 9.94452
R21 R2R_20k_0.B1.n1 R2R_20k_0.B1.t5 2.36193
R22 R2R_20k_0.B1.n1 R2R_20k_0.B1.t0 2.36193
R23 R2R_20k_0.B1.n4 R2R_20k_0.B1.n3 1.83465
R24 R2R_20k_0.B1.n4 R2R_20k_0.B1.n2 1.82789
R25 R2R_20k_0.B1.n0 R2R_20k_0.B1.t1 1.73144
R26 R2R_20k_0.B1.n0 R2R_20k_0.B1.t2 1.73144
R27 R2R_20k_0.B1.n5 R2R_20k_0.B1 0.80378
R28 R2R_20k_0.B1 R2R_20k_0.B1.n4 0.0623812
R29 R2R_20k_0.B1 R2R_20k_0.B1.n5 0.06175
R30 V_REF.n27 V_REF.n21 6832.14
R31 V_REF.n17 V_REF.n16 6832.14
R32 V_REF.n37 V_REF.n15 6832.14
R33 V_REF.n11 V_REF.n10 6832.14
R34 V_REF.n47 V_REF.n9 6832.14
R35 V_REF.n48 V_REF.n5 6832.14
R36 V_REF.n3 V_REF.n2 6710.8
R37 V_REF.n27 V_REF.n26 749.662
R38 V_REF.n28 V_REF.n27 729.207
R39 V_REF.n28 V_REF.n16 729.207
R40 V_REF.n36 V_REF.n16 729.207
R41 V_REF.n37 V_REF.n36 729.207
R42 V_REF.n38 V_REF.n37 729.207
R43 V_REF.n38 V_REF.n10 729.207
R44 V_REF.n46 V_REF.n10 729.207
R45 V_REF.n47 V_REF.n46 729.207
R46 V_REF.n49 V_REF.n47 729.207
R47 V_REF.n49 V_REF.n48 729.207
R48 V_REF.n48 V_REF.n4 729.207
R49 V_REF.n25 V_REF.n21 729.207
R50 V_REF.n29 V_REF.n21 729.207
R51 V_REF.n29 V_REF.n17 729.207
R52 V_REF.n35 V_REF.n17 729.207
R53 V_REF.n35 V_REF.n15 729.207
R54 V_REF.n39 V_REF.n15 729.207
R55 V_REF.n39 V_REF.n11 729.207
R56 V_REF.n45 V_REF.n11 729.207
R57 V_REF.n45 V_REF.n9 729.207
R58 V_REF.n50 V_REF.n9 729.207
R59 V_REF.n50 V_REF.n5 729.207
R60 V_REF.n57 V_REF.n5 729.207
R61 V_REF.n58 V_REF.n3 692.532
R62 V_REF.n57 V_REF.n2 672.077
R63 V_REF.n59 V_REF.n2 668.277
R64 V_REF.n4 V_REF.n3 668.277
R65 V_REF.t30 V_REF.t16 108.674
R66 V_REF.t26 V_REF.t20 108.674
R67 V_REF.t18 V_REF.t10 108.674
R68 V_REF.t44 V_REF.t2 108.674
R69 V_REF.t34 V_REF.t4 108.674
R70 V_REF.t24 V_REF.t38 108.674
R71 V_REF.t22 V_REF.t40 108.15
R72 V_REF.t46 V_REF.t28 40.3066
R73 V_REF.t46 V_REF.t30 40.3066
R74 V_REF.t32 V_REF.t16 40.3066
R75 V_REF.t32 V_REF.t26 40.3066
R76 V_REF.t8 V_REF.t20 40.3066
R77 V_REF.t8 V_REF.t18 40.3066
R78 V_REF.t36 V_REF.t10 40.3066
R79 V_REF.t36 V_REF.t44 40.3066
R80 V_REF.t0 V_REF.t2 40.3066
R81 V_REF.t0 V_REF.t34 40.3066
R82 V_REF.t12 V_REF.t4 40.3066
R83 V_REF.t12 V_REF.t24 40.3066
R84 V_REF.t42 V_REF.t38 40.3066
R85 V_REF.t40 V_REF.t42 40.3066
R86 V_REF.t6 V_REF.t22 40.3066
R87 V_REF.t6 V_REF.t14 40.3066
R88 V_REF.n25 V_REF.n24 21.5894
R89 V_REF.n30 V_REF.n29 21.5894
R90 V_REF.n35 V_REF.n34 21.5894
R91 V_REF.n40 V_REF.n39 21.5894
R92 V_REF.n45 V_REF.n44 21.5894
R93 V_REF.n51 V_REF.n50 21.5894
R94 V_REF.n57 V_REF.n56 21.5894
R95 V_REF.n60 V_REF.n59 21.5894
R96 V_REF.t42 V_REF.n4 20.5561
R97 V_REF.t12 V_REF.n49 20.5561
R98 V_REF.n46 V_REF.t0 20.5561
R99 V_REF.t36 V_REF.n38 20.5561
R100 V_REF.n36 V_REF.t8 20.5561
R101 V_REF.t32 V_REF.n28 20.5561
R102 V_REF.n29 V_REF.t32 20.5561
R103 V_REF.t8 V_REF.n35 20.5561
R104 V_REF.n39 V_REF.t36 20.5561
R105 V_REF.t0 V_REF.n45 20.5561
R106 V_REF.n50 V_REF.t12 20.5561
R107 V_REF.t42 V_REF.n57 20.5561
R108 V_REF.n59 V_REF.n58 20.4551
R109 V_REF.n26 V_REF.n25 20.4551
R110 V_REF.n55 V_REF.t41 18.9603
R111 V_REF.n52 V_REF.t25 18.9603
R112 V_REF.n43 V_REF.t35 18.9603
R113 V_REF.n41 V_REF.t45 18.9603
R114 V_REF.n33 V_REF.t19 18.9603
R115 V_REF.n31 V_REF.t27 18.9603
R116 V_REF.n23 V_REF.t31 18.9603
R117 V_REF.n61 V_REF.t15 18.9548
R118 V_REF.n24 V_REF.n22 17.2568
R119 V_REF.n53 V_REF.n6 17.2293
R120 V_REF.n8 V_REF.n7 17.2293
R121 V_REF.n42 V_REF.n12 17.2293
R122 V_REF.n14 V_REF.n13 17.2293
R123 V_REF.n32 V_REF.n18 17.2293
R124 V_REF.n20 V_REF.n19 17.2293
R125 V_REF.n1 V_REF.n0 17.2293
R126 V_REF.n6 V_REF.t39 1.73144
R127 V_REF.n6 V_REF.t43 1.73144
R128 V_REF.n7 V_REF.t5 1.73144
R129 V_REF.n7 V_REF.t13 1.73144
R130 V_REF.n12 V_REF.t3 1.73144
R131 V_REF.n12 V_REF.t1 1.73144
R132 V_REF.n13 V_REF.t11 1.73144
R133 V_REF.n13 V_REF.t37 1.73144
R134 V_REF.n18 V_REF.t21 1.73144
R135 V_REF.n18 V_REF.t9 1.73144
R136 V_REF.n19 V_REF.t17 1.73144
R137 V_REF.n19 V_REF.t33 1.73144
R138 V_REF.n22 V_REF.t29 1.73144
R139 V_REF.n22 V_REF.t47 1.73144
R140 V_REF.n0 V_REF.t23 1.73144
R141 V_REF.n0 V_REF.t7 1.73144
R142 V_REF V_REF.n20 0.0918194
R143 V_REF.n32 V_REF 0.0918194
R144 V_REF V_REF.n14 0.0918194
R145 V_REF.n42 V_REF 0.0918194
R146 V_REF V_REF.n8 0.0918194
R147 V_REF.n53 V_REF 0.0918194
R148 V_REF V_REF.n1 0.0906243
R149 V_REF.n24 V_REF.n23 0.0827917
R150 V_REF.n31 V_REF.n30 0.0827917
R151 V_REF.n34 V_REF.n33 0.0827917
R152 V_REF.n41 V_REF.n40 0.0827917
R153 V_REF.n44 V_REF.n43 0.0827917
R154 V_REF.n52 V_REF.n51 0.0827917
R155 V_REF.n56 V_REF.n55 0.0827917
R156 V_REF.n61 V_REF.n60 0.0821909
R157 V_REF.n23 V_REF 0.0570972
R158 V_REF V_REF.n31 0.0570972
R159 V_REF.n33 V_REF 0.0570972
R160 V_REF V_REF.n41 0.0570972
R161 V_REF.n43 V_REF 0.0570972
R162 V_REF V_REF.n52 0.0570972
R163 V_REF V_REF.n61 0.0564753
R164 V_REF.n58 V_REF.t6 0.0517139
R165 V_REF.n26 V_REF.t46 0.0517139
R166 V_REF.n55 V_REF.n54 0.0362639
R167 V_REF.n30 V_REF.n20 0.0279306
R168 V_REF.n34 V_REF.n32 0.0279306
R169 V_REF.n40 V_REF.n14 0.0279306
R170 V_REF.n44 V_REF.n42 0.0279306
R171 V_REF.n51 V_REF.n8 0.0279306
R172 V_REF.n56 V_REF.n53 0.0279306
R173 V_REF.n60 V_REF.n1 0.027779
R174 V_REF.n54 V_REF 0.0213333
R175 V_REF.n54 V_REF 0.0212182
R176 V_COM.n71 V_COM.n3 284216
R177 V_COM.n72 V_COM.n2 12851.4
R178 V_COM.n26 V_COM.n2 12851.4
R179 V_COM.n27 V_COM.n2 6425.68
R180 V_COM.n11 V_COM.n10 5486.31
R181 V_COM.n52 V_COM.n15 5486.31
R182 V_COM.n17 V_COM.n16 5486.31
R183 V_COM.n42 V_COM.n21 5486.31
R184 V_COM.n23 V_COM.n22 5486.31
R185 V_COM.n62 V_COM.n9 5486.31
R186 V_COM.n5 V_COM.n4 5481.7
R187 V_COM.n33 V_COM.n22 1285.69
R188 V_COM.n41 V_COM.n22 1221.74
R189 V_COM.n42 V_COM.n41 1221.74
R190 V_COM.n43 V_COM.n42 1221.74
R191 V_COM.n43 V_COM.n16 1221.74
R192 V_COM.n51 V_COM.n16 1221.74
R193 V_COM.n52 V_COM.n51 1221.74
R194 V_COM.n53 V_COM.n52 1221.74
R195 V_COM.n53 V_COM.n10 1221.74
R196 V_COM.n61 V_COM.n10 1221.74
R197 V_COM.n62 V_COM.n61 1221.74
R198 V_COM.n63 V_COM.n62 1221.74
R199 V_COM.n34 V_COM.n23 1221.74
R200 V_COM.n40 V_COM.n23 1221.74
R201 V_COM.n40 V_COM.n21 1221.74
R202 V_COM.n44 V_COM.n21 1221.74
R203 V_COM.n44 V_COM.n17 1221.74
R204 V_COM.n50 V_COM.n17 1221.74
R205 V_COM.n50 V_COM.n15 1221.74
R206 V_COM.n54 V_COM.n15 1221.74
R207 V_COM.n54 V_COM.n11 1221.74
R208 V_COM.n60 V_COM.n11 1221.74
R209 V_COM.n60 V_COM.n9 1221.74
R210 V_COM.n64 V_COM.n9 1221.74
R211 V_COM.n70 V_COM.n4 1183.61
R212 V_COM.n69 V_COM.n5 1126.02
R213 V_COM.n63 V_COM.n4 1126.02
R214 V_COM.n64 V_COM.n5 1119.66
R215 V_COM.t2 V_COM.t36 211.852
R216 V_COM.t76 V_COM.t67 211.852
R217 V_COM.t25 V_COM.t70 211.766
R218 V_COM.t5 V_COM.t38 211.766
R219 V_COM.t66 V_COM.t79 211.766
R220 V_COM.t41 V_COM.t4 211.766
R221 V_COM.t42 V_COM.t3 211.766
R222 V_COM.t69 V_COM.t30 211.766
R223 V_COM.t6 V_COM.t65 201.81
R224 V_COM.t65 V_COM.t74 183.71
R225 V_COM.t19 V_COM.t69 165.612
R226 V_COM.t42 V_COM.t23 147.512
R227 V_COM.t53 V_COM.t9 143.046
R228 V_COM.t34 V_COM.t39 142.987
R229 V_COM.t0 V_COM.t26 142.987
R230 V_COM.t31 V_COM.t44 142.987
R231 V_COM.t55 V_COM.t17 142.987
R232 V_COM.t59 V_COM.t61 142.987
R233 V_COM.t70 V_COM.n3 138.463
R234 V_COM.t48 V_COM.t50 136.653
R235 V_COM.t51 V_COM.t5 134.843
R236 V_COM.t28 V_COM.t46 133.032
R237 V_COM.t63 V_COM.t2 117.198
R238 V_COM.t11 V_COM.t58 116.79
R239 V_COM.t13 V_COM.t73 114.933
R240 V_COM.t8 V_COM.t21 113.123
R241 V_COM.t4 V_COM.t15 111.312
R242 V_COM.t15 V_COM.t37 100.453
R243 V_COM.t21 V_COM.t66 98.643
R244 V_COM.t13 V_COM.t43 96.8331
R245 V_COM.t67 V_COM.t11 95.0622
R246 V_COM.n71 V_COM.t76 94.1569
R247 V_COM.n72 V_COM.n71 87.8237
R248 V_COM.t47 V_COM.t63 82.3534
R249 V_COM.t28 V_COM.t33 78.7335
R250 V_COM.t57 V_COM.t51 76.9236
R251 V_COM.t79 V_COM.t48 75.1136
R252 V_COM.t34 V_COM.t57 66.0639
R253 V_COM.n65 V_COM.n64 66.0338
R254 V_COM.n60 V_COM.n59 66.0338
R255 V_COM.n55 V_COM.n54 66.0338
R256 V_COM.n50 V_COM.n49 66.0338
R257 V_COM.n45 V_COM.n44 66.0338
R258 V_COM.n40 V_COM.n39 66.0338
R259 V_COM.n35 V_COM.n34 66.0338
R260 V_COM.n69 V_COM.n68 66.0338
R261 V_COM.n64 V_COM.t59 65.0005
R262 V_COM.t13 V_COM.n60 65.0005
R263 V_COM.n54 V_COM.t28 65.0005
R264 V_COM.t55 V_COM.n50 65.0005
R265 V_COM.n44 V_COM.t31 65.0005
R266 V_COM.t0 V_COM.n40 65.0005
R267 V_COM.n41 V_COM.t0 65.0005
R268 V_COM.t31 V_COM.n43 65.0005
R269 V_COM.n51 V_COM.t55 65.0005
R270 V_COM.t28 V_COM.n53 65.0005
R271 V_COM.n61 V_COM.t13 65.0005
R272 V_COM.t59 V_COM.n63 65.0005
R273 V_COM.t23 V_COM.t33 64.2539
R274 V_COM.n70 V_COM.n69 63.9526
R275 V_COM.n34 V_COM.n33 63.9526
R276 V_COM.t44 V_COM.t41 62.4439
R277 V_COM.t59 V_COM.t47 60.634
R278 V_COM.t43 V_COM.t19 46.1543
R279 V_COM.n26 V_COM.n3 43.4507
R280 V_COM.t36 V_COM.t9 42.5519
R281 V_COM.t55 V_COM.t37 42.5344
R282 V_COM.t38 V_COM.t26 38.9145
R283 V_COM.t0 V_COM.t8 29.8648
R284 V_COM.t74 V_COM.t73 28.0548
R285 V_COM.t58 V_COM.t53 26.2556
R286 V_COM.t3 V_COM.t17 26.2448
R287 V_COM.n1 V_COM.t78 21.5736
R288 V_COM.n29 V_COM.t72 21.5736
R289 V_COM.n31 V_COM.t71 21.4809
R290 V_COM.n74 V_COM.t68 21.4809
R291 V_COM.n74 V_COM.t77 21.4809
R292 V_COM.n30 V_COM.n26 17.6313
R293 V_COM.n73 V_COM.n72 17.497
R294 V_COM.n36 V_COM.t52 14.2264
R295 V_COM.n38 V_COM.t22 14.2264
R296 V_COM.n46 V_COM.t45 14.2264
R297 V_COM.n48 V_COM.t18 14.2264
R298 V_COM.n56 V_COM.t7 14.2264
R299 V_COM.n58 V_COM.t20 14.2264
R300 V_COM.n66 V_COM.t64 14.2264
R301 V_COM.n0 V_COM.t12 14.221
R302 V_COM.n32 V_COM.n25 11.865
R303 V_COM.n37 V_COM.n24 11.865
R304 V_COM.n20 V_COM.n19 11.865
R305 V_COM.n47 V_COM.n18 11.865
R306 V_COM.n14 V_COM.n13 11.865
R307 V_COM.n57 V_COM.n12 11.865
R308 V_COM.n8 V_COM.n7 11.865
R309 V_COM.n67 V_COM.n6 11.8595
R310 V_COM.t46 V_COM.t6 9.95525
R311 V_COM.t30 V_COM.t61 8.1453
R312 V_COM.n28 V_COM.n27 6.39772
R313 V_COM.t31 V_COM.t50 6.33534
R314 V_COM.n27 V_COM.t42 6.29082
R315 V_COM.n29 V_COM.n28 4.66286
R316 V_COM.n28 V_COM.n1 4.19278
R317 V_COM.t39 V_COM.t25 2.71543
R318 V_COM.n25 V_COM.t40 2.36193
R319 V_COM.n25 V_COM.t35 2.36193
R320 V_COM.n24 V_COM.t27 2.36193
R321 V_COM.n24 V_COM.t1 2.36193
R322 V_COM.n19 V_COM.t49 2.36193
R323 V_COM.n19 V_COM.t32 2.36193
R324 V_COM.n18 V_COM.t16 2.36193
R325 V_COM.n18 V_COM.t56 2.36193
R326 V_COM.n13 V_COM.t24 2.36193
R327 V_COM.n13 V_COM.t29 2.36193
R328 V_COM.n12 V_COM.t75 2.36193
R329 V_COM.n12 V_COM.t14 2.36193
R330 V_COM.n7 V_COM.t62 2.36193
R331 V_COM.n7 V_COM.t60 2.36193
R332 V_COM.n6 V_COM.t10 2.36193
R333 V_COM.n6 V_COM.t54 2.36193
R334 V_COM.n30 V_COM.n29 2.21144
R335 V_COM.n32 V_COM.n31 1.50825
R336 V_COM.n31 V_COM.n30 1.30323
R337 V_COM.n33 V_COM.t34 0.525207
R338 V_COM.t53 V_COM.n70 0.525207
R339 V_COM.n73 V_COM.n1 0.402286
R340 V_COM.n74 V_COM.n73 0.358757
R341 V_COM.n76 V_COM 0.268288
R342 V_COM.n76 V_COM.n75 0.17164
R343 V_COM.n37 V_COM 0.136347
R344 V_COM V_COM.n20 0.136347
R345 V_COM.n47 V_COM 0.136347
R346 V_COM V_COM.n14 0.136347
R347 V_COM.n57 V_COM 0.136347
R348 V_COM V_COM.n8 0.136347
R349 V_COM.n67 V_COM 0.135314
R350 V_COM.n36 V_COM.n35 0.122917
R351 V_COM.n39 V_COM.n38 0.122917
R352 V_COM.n46 V_COM.n45 0.122917
R353 V_COM.n49 V_COM.n48 0.122917
R354 V_COM.n56 V_COM.n55 0.122917
R355 V_COM.n59 V_COM.n58 0.122917
R356 V_COM.n66 V_COM.n65 0.122917
R357 V_COM.n68 V_COM.n0 0.122917
R358 V_COM.n75 V_COM.n74 0.120277
R359 V_COM V_COM.n36 0.0846942
R360 V_COM.n38 V_COM 0.0846942
R361 V_COM V_COM.n46 0.0846942
R362 V_COM.n48 V_COM 0.0846942
R363 V_COM V_COM.n56 0.0846942
R364 V_COM.n58 V_COM 0.0846942
R365 V_COM V_COM.n66 0.0846942
R366 V_COM V_COM.n0 0.0846942
R367 V_COM.n75 V_COM 0.0578347
R368 V_COM.n35 V_COM.n32 0.0413058
R369 V_COM.n39 V_COM.n37 0.0413058
R370 V_COM.n45 V_COM.n20 0.0413058
R371 V_COM.n49 V_COM.n47 0.0413058
R372 V_COM.n55 V_COM.n14 0.0413058
R373 V_COM.n59 V_COM.n57 0.0413058
R374 V_COM.n65 V_COM.n8 0.0413058
R375 V_COM.n68 V_COM.n67 0.0413058
R376 V_COM V_COM.n76 0.0247769
R377 D0.n5 D0.t1 963.587
R378 D0.n0 D0.t3 963.587
R379 D0.n1 D0.t0 963.587
R380 D0.n2 D0.t2 515.91
R381 D0.n3 D0.t5 515.91
R382 D0.n4 D0.t4 515.91
R383 D0.n4 D0.n3 59.4829
R384 D0.n3 D0.n2 59.4829
R385 D0.n3 D0.n0 9.54099
R386 D0.n5 D0.n4 9.54099
R387 D0.n2 D0.n1 9.54099
R388 D0 D0.n6 7.34316
R389 D0 D0.n0 0.063
R390 D0.n6 D0.n0 0.0506312
R391 D0.n6 D0.n5 0.050027
R392 D0.n1 D0 0.03675
R393 R2R_20k_0.B0.n5 R2R_20k_0.B0.t0 21.7118
R394 R2R_20k_0.B0.n3 R2R_20k_0.B0.t5 20.8848
R395 R2R_20k_0.B0.n2 R2R_20k_0.B0.n0 19.1576
R396 R2R_20k_0.B0.n3 R2R_20k_0.B0.t2 12.3059
R397 R2R_20k_0.B0.n2 R2R_20k_0.B0.n1 9.94452
R398 R2R_20k_0.B0.n1 R2R_20k_0.B0.t1 2.36193
R399 R2R_20k_0.B0.n1 R2R_20k_0.B0.t3 2.36193
R400 R2R_20k_0.B0.n4 R2R_20k_0.B0.n3 1.83828
R401 R2R_20k_0.B0.n4 R2R_20k_0.B0.n2 1.82473
R402 R2R_20k_0.B0.n0 R2R_20k_0.B0.t4 1.73144
R403 R2R_20k_0.B0.n0 R2R_20k_0.B0.t6 1.73144
R404 R2R_20k_0.B0.n5 R2R_20k_0.B0 0.827639
R405 R2R_20k_0.B0 R2R_20k_0.B0.n4 0.0623812
R406 R2R_20k_0.B0 R2R_20k_0.B0.n5 0.061125
R407 D5.n5 D5.t1 963.587
R408 D5.n0 D5.t0 963.587
R409 D5.n1 D5.t3 963.587
R410 D5.n2 D5.t5 515.91
R411 D5.n3 D5.t2 515.91
R412 D5.n4 D5.t4 515.91
R413 D5.n4 D5.n3 59.4829
R414 D5.n3 D5.n2 59.4829
R415 D5.n3 D5.n0 9.54099
R416 D5.n5 D5.n4 9.54099
R417 D5.n2 D5.n1 9.54099
R418 D5 D5.n6 7.5689
R419 D5 D5.n0 0.063
R420 D5.n6 D5.n5 0.0575721
R421 D5.n6 D5.n0 0.0431329
R422 D5.n1 D5 0.03675
R423 R2R_20k_0.B5.n5 R2R_20k_0.B5.t6 21.7179
R424 R2R_20k_0.B5.n3 R2R_20k_0.B5.t4 20.8848
R425 R2R_20k_0.B5.n2 R2R_20k_0.B5.n0 19.1576
R426 R2R_20k_0.B5.n3 R2R_20k_0.B5.t1 12.3059
R427 R2R_20k_0.B5.n2 R2R_20k_0.B5.n1 9.94452
R428 R2R_20k_0.B5.n1 R2R_20k_0.B5.t2 2.36193
R429 R2R_20k_0.B5.n1 R2R_20k_0.B5.t0 2.36193
R430 R2R_20k_0.B5.n4 R2R_20k_0.B5.n3 1.83828
R431 R2R_20k_0.B5.n4 R2R_20k_0.B5.n2 1.82473
R432 R2R_20k_0.B5.n0 R2R_20k_0.B5.t5 1.73144
R433 R2R_20k_0.B5.n0 R2R_20k_0.B5.t3 1.73144
R434 R2R_20k_0.B5.n5 R2R_20k_0.B5 0.703804
R435 R2R_20k_0.B5 R2R_20k_0.B5.n4 0.0623812
R436 R2R_20k_0.B5 R2R_20k_0.B5.n5 0.0623812
R437 D7.n5 D7.t3 963.587
R438 D7.n0 D7.t2 963.587
R439 D7.n1 D7.t4 963.587
R440 D7.n2 D7.t1 515.91
R441 D7.n3 D7.t5 515.91
R442 D7.n4 D7.t0 515.91
R443 D7.n4 D7.n3 59.4829
R444 D7.n3 D7.n2 59.4829
R445 D7.n3 D7.n0 9.54099
R446 D7.n5 D7.n4 9.54099
R447 D7.n2 D7.n1 9.54099
R448 D7 D7.n6 7.5689
R449 D7 D7.n0 0.063
R450 D7.n6 D7.n5 0.0600721
R451 D7.n6 D7.n0 0.0406329
R452 D7.n1 D7 0.03675
R453 R2R_20k_0.B7.n5 R2R_20k_0.B7.t0 21.7166
R454 R2R_20k_0.B7.n0 R2R_20k_0.B7.t5 20.8848
R455 R2R_20k_0.B7.n3 R2R_20k_0.B7.n1 19.1576
R456 R2R_20k_0.B7.n0 R2R_20k_0.B7.t3 12.3059
R457 R2R_20k_0.B7.n3 R2R_20k_0.B7.n2 9.94452
R458 R2R_20k_0.B7.n2 R2R_20k_0.B7.t1 2.36193
R459 R2R_20k_0.B7.n2 R2R_20k_0.B7.t2 2.36193
R460 R2R_20k_0.B7.n4 R2R_20k_0.B7.n0 1.73397
R461 R2R_20k_0.B7.n1 R2R_20k_0.B7.t6 1.73144
R462 R2R_20k_0.B7.n1 R2R_20k_0.B7.t4 1.73144
R463 R2R_20k_0.B7 R2R_20k_0.B7.n3 1.72397
R464 R2R_20k_0.B7.n5 R2R_20k_0.B7.n4 0.6905
R465 R2R_20k_0.B7.n4 R2R_20k_0.B7 0.11175
R466 R2R_20k_0.B7 R2R_20k_0.B7.n5 0.063
R467 R2R_20k_0.B6.n5 R2R_20k_0.B6.t5 21.7164
R468 R2R_20k_0.B6.n0 R2R_20k_0.B6.t2 20.8848
R469 R2R_20k_0.B6.n3 R2R_20k_0.B6.n1 19.1576
R470 R2R_20k_0.B6.n0 R2R_20k_0.B6.t3 12.3059
R471 R2R_20k_0.B6.n3 R2R_20k_0.B6.n2 9.94452
R472 R2R_20k_0.B6.n2 R2R_20k_0.B6.t0 2.36193
R473 R2R_20k_0.B6.n2 R2R_20k_0.B6.t1 2.36193
R474 R2R_20k_0.B6.n4 R2R_20k_0.B6.n0 1.78272
R475 R2R_20k_0.B6.n1 R2R_20k_0.B6.t6 1.73144
R476 R2R_20k_0.B6.n1 R2R_20k_0.B6.t4 1.73144
R477 R2R_20k_0.B6 R2R_20k_0.B6.n3 1.72397
R478 R2R_20k_0.B6.n5 R2R_20k_0.B6.n4 0.686502
R479 R2R_20k_0.B6.n4 R2R_20k_0.B6 0.063
R480 R2R_20k_0.B6 R2R_20k_0.B6.n5 0.0617624
R481 D4.n5 D4.t0 963.587
R482 D4.n0 D4.t1 963.587
R483 D4.n1 D4.t5 963.587
R484 D4.n2 D4.t2 515.91
R485 D4.n3 D4.t3 515.91
R486 D4.n4 D4.t4 515.91
R487 D4.n4 D4.n3 59.4829
R488 D4.n3 D4.n2 59.4829
R489 D4.n3 D4.n0 9.54099
R490 D4.n5 D4.n4 9.54099
R491 D4.n2 D4.n1 9.54099
R492 D4 D4.n6 7.56792
R493 D4 D4.n0 0.063
R494 D4.n6 D4.n5 0.0571483
R495 D4.n6 D4.n0 0.04355
R496 D4.n1 D4 0.03675
R497 R2R_20k_0.B4.n5 R2R_20k_0.B4.t0 21.716
R498 R2R_20k_0.B4.n0 R2R_20k_0.B4.t6 20.8848
R499 R2R_20k_0.B4.n3 R2R_20k_0.B4.n1 19.1576
R500 R2R_20k_0.B4.n0 R2R_20k_0.B4.t1 12.3059
R501 R2R_20k_0.B4.n3 R2R_20k_0.B4.n2 9.94452
R502 R2R_20k_0.B4.n2 R2R_20k_0.B4.t2 2.36193
R503 R2R_20k_0.B4.n2 R2R_20k_0.B4.t3 2.36193
R504 R2R_20k_0.B4.n4 R2R_20k_0.B4.n0 1.78397
R505 R2R_20k_0.B4.n1 R2R_20k_0.B4.t5 1.73144
R506 R2R_20k_0.B4.n1 R2R_20k_0.B4.t4 1.73144
R507 R2R_20k_0.B4 R2R_20k_0.B4.n3 1.72397
R508 R2R_20k_0.B4.n5 R2R_20k_0.B4.n4 0.734858
R509 R2R_20k_0.B4 R2R_20k_0.B4.n5 0.063
R510 R2R_20k_0.B4.n4 R2R_20k_0.B4 0.06175
R511 D2.n5 D2.t4 963.587
R512 D2.n0 D2.t3 963.587
R513 D2.n1 D2.t0 963.587
R514 D2.n2 D2.t2 515.91
R515 D2.n3 D2.t5 515.91
R516 D2.n4 D2.t1 515.91
R517 D2.n4 D2.n3 59.4829
R518 D2.n3 D2.n2 59.4829
R519 D2.n3 D2.n0 9.54099
R520 D2.n5 D2.n4 9.54099
R521 D2.n2 D2.n1 9.54099
R522 D2 D2.n6 7.5684
R523 D2 D2.n0 0.063
R524 D2.n6 D2.n5 0.0592352
R525 D2.n6 D2.n0 0.0414665
R526 D2.n1 D2 0.03675
R527 R2R_20k_0.B2.n5 R2R_20k_0.B2.t6 21.7063
R528 R2R_20k_0.B2.n0 R2R_20k_0.B2.t3 20.8848
R529 R2R_20k_0.B2.n3 R2R_20k_0.B2.n1 19.1576
R530 R2R_20k_0.B2.n0 R2R_20k_0.B2.t2 12.3059
R531 R2R_20k_0.B2.n3 R2R_20k_0.B2.n2 9.94452
R532 R2R_20k_0.B2.n2 R2R_20k_0.B2.t0 2.36193
R533 R2R_20k_0.B2.n2 R2R_20k_0.B2.t1 2.36193
R534 R2R_20k_0.B2.n4 R2R_20k_0.B2.n0 1.78209
R535 R2R_20k_0.B2.n1 R2R_20k_0.B2.t4 1.73144
R536 R2R_20k_0.B2.n1 R2R_20k_0.B2.t5 1.73144
R537 R2R_20k_0.B2 R2R_20k_0.B2.n3 1.72397
R538 R2R_20k_0.B2.n5 R2R_20k_0.B2.n4 0.779793
R539 R2R_20k_0.B2.n4 R2R_20k_0.B2 0.063625
R540 R2R_20k_0.B2 R2R_20k_0.B2.n5 0.063625
R541 D6.n5 D6.t1 963.587
R542 D6.n0 D6.t2 963.587
R543 D6.n1 D6.t0 963.587
R544 D6.n2 D6.t4 515.91
R545 D6.n3 D6.t5 515.91
R546 D6.n4 D6.t3 515.91
R547 D6.n4 D6.n3 59.4829
R548 D6.n3 D6.n2 59.4829
R549 D6.n3 D6.n0 9.54099
R550 D6.n5 D6.n4 9.54099
R551 D6.n2 D6.n1 9.54099
R552 D6 D6.n6 7.57046
R553 D6 D6.n0 0.063
R554 D6.n6 D6.n5 0.0575824
R555 D6.n6 D6.n0 0.0431317
R556 D6.n1 D6 0.03675
R557 D3.n5 D3.t1 963.587
R558 D3.n0 D3.t4 963.587
R559 D3.n1 D3.t5 963.587
R560 D3.n2 D3.t2 515.91
R561 D3.n3 D3.t3 515.91
R562 D3.n4 D3.t0 515.91
R563 D3.n4 D3.n3 59.4829
R564 D3.n3 D3.n2 59.4829
R565 D3.n3 D3.n0 9.54099
R566 D3.n5 D3.n4 9.54099
R567 D3.n2 D3.n1 9.54099
R568 D3 D3.n6 7.5684
R569 D3 D3.n0 0.063
R570 D3.n6 D3.n5 0.0592352
R571 D3.n6 D3.n0 0.0414665
R572 D3.n1 D3 0.03675
R573 R2R_20k_0.B3.n5 R2R_20k_0.B3.t0 21.71
R574 R2R_20k_0.B3.n3 R2R_20k_0.B3.t6 20.8848
R575 R2R_20k_0.B3.n2 R2R_20k_0.B3.n0 19.1576
R576 R2R_20k_0.B3.n3 R2R_20k_0.B3.t3 12.3059
R577 R2R_20k_0.B3.n2 R2R_20k_0.B3.n1 9.94452
R578 R2R_20k_0.B3.n1 R2R_20k_0.B3.t1 2.36193
R579 R2R_20k_0.B3.n1 R2R_20k_0.B3.t2 2.36193
R580 R2R_20k_0.B3.n4 R2R_20k_0.B3.n3 1.83828
R581 R2R_20k_0.B3.n4 R2R_20k_0.B3.n2 1.82789
R582 R2R_20k_0.B3.n0 R2R_20k_0.B3.t5 1.73144
R583 R2R_20k_0.B3.n0 R2R_20k_0.B3.t4 1.73144
R584 R2R_20k_0.B3.n5 R2R_20k_0.B3 0.758109
R585 R2R_20k_0.B3 R2R_20k_0.B3.n5 0.063
R586 R2R_20k_0.B3 R2R_20k_0.B3.n4 0.0617745
R587 V_out.n0 V_out.t1 21.4809
R588 V_out.n0 V_out.t0 21.4809
R589 V_out V_out.n1 0.395602
R590 V_out.n1 V_out 0.0403649
R591 V_out.n1 V_out.n0 0.035973
C0 a_n798_n2638# a_n330_n2638# 0.296492f
C1 V_REF D2 2.31853f
C2 R2R_20k_0.B0 D2 3.08e-20
C3 D1 R2R_20k_0.B1 4.247f
C4 R2R_20k_0.B3 R2R_20k_0.B4 0.717628f
C5 a_2478_n2638# a_1776_n2638# 3.82e-20
C6 D0 R2R_20k_0.B1 4.65e-19
C7 a_2946_n838# a_2244_n838# 0.128514f
C8 m4_n961_5637# V_REF 0.134033f
C9 D6 V_REF 2.31839f
C10 a_1074_n2638# a_372_n2638# 3.02e-19
C11 a_3648_n838# R2R_20k_0.B6 0.335561f
C12 R2R_20k_0.B7 V_REF 4.92015f
C13 D0 a_n564_n838# 0.001264f
C14 a_2244_n838# R2R_20k_0.B4 0.376318f
C15 D3 D2 0.115681f
C16 R2R_20k_0.B1 R2R_20k_0.B3 1.96e-19
C17 a_1074_n2638# a_840_n838# 0.402638f
C18 V_out R2R_20k_0.B6 0.466537f
C19 D4 R2R_20k_0.B4 4.25967f
C20 D1 V_REF 2.31922f
C21 D1 R2R_20k_0.B0 0.017497f
C22 D6 D5 0.115763f
C23 a_3648_n838# R2R_20k_0.B5 0.300007f
C24 a_2244_n838# R2R_20k_0.B3 0.298919f
C25 R2R_20k_0.B3 a_840_n838# 5.1e-20
C26 D0 V_REF 2.39944f
C27 R2R_20k_0.B1 a_372_n2638# 0.002521f
C28 D0 R2R_20k_0.B0 4.40085f
C29 D4 R2R_20k_0.B3 0.016236f
C30 a_3648_n838# a_4584_n2638# 0.299255f
C31 V_REF R2R_20k_0.B4 5.8023f
C32 D7 V_out 0.007847f
C33 V_out R2R_20k_0.B5 1.33e-19
C34 a_3180_n2638# R2R_20k_0.B5 0.002521f
C35 D6 R2R_20k_0.B6 4.24985f
C36 a_2946_n838# D5 0.001396f
C37 a_n564_n838# R2R_20k_0.B1 2.75e-21
C38 R2R_20k_0.B2 D2 4.25162f
C39 R2R_20k_0.B7 R2R_20k_0.B6 0.664267f
C40 a_4584_n2638# V_out 0.00699f
C41 R2R_20k_0.B1 a_840_n838# 0.299419f
C42 a_n564_n838# a_372_n2638# 0.299243f
C43 V_REF R2R_20k_0.B3 5.80222f
C44 a_840_n838# a_372_n2638# 1.19e-20
C45 R2R_20k_0.B3 a_1542_n838# 0.404376f
C46 D5 R2R_20k_0.B4 0.016236f
C47 D7 D6 0.115762f
C48 D6 R2R_20k_0.B5 0.016236f
C49 D4 a_2244_n838# 0.001304f
C50 R2R_20k_0.B7 D7 4.2488f
C51 R2R_20k_0.B1 V_REF 5.80224f
C52 R2R_20k_0.B0 R2R_20k_0.B1 0.741772f
C53 R2R_20k_0.B1 a_1542_n838# 1.78e-20
C54 D3 R2R_20k_0.B4 1.99e-19
C55 a_1542_n838# a_372_n2638# 2.46e-21
C56 R2R_20k_0.B7 a_4584_n2638# 0.006187f
C57 a_3180_n2638# a_1776_n2638# 6.25e-21
C58 a_2946_n838# R2R_20k_0.B5 0.35707f
C59 a_n564_n838# R2R_20k_0.B0 0.4593f
C60 a_2244_n838# a_1542_n838# 0.127701f
C61 R2R_20k_0.B2 D1 1.99e-19
C62 D3 R2R_20k_0.B3 4.25169f
C63 a_2478_n2638# R2R_20k_0.B4 0.002521f
C64 a_1542_n838# a_840_n838# 0.131021f
C65 D4 V_REF 2.31642f
C66 a_3882_n2638# R2R_20k_0.B6 0.002521f
C67 R2R_20k_0.B5 R2R_20k_0.B4 0.713568f
C68 R2R_20k_0.B2 D0 1.33e-20
C69 R2R_20k_0.B2 R2R_20k_0.B4 9.84e-21
C70 R2R_20k_0.B2 a_1074_n2638# 0.002521f
C71 R2R_20k_0.B0 V_REF 5.80799f
C72 D4 D5 0.115764f
C73 R2R_20k_0.B5 R2R_20k_0.B3 9.39e-20
C74 a_3648_n838# V_out 0.008425f
C75 a_2946_n838# a_1776_n2638# 1.26e-21
C76 R2R_20k_0.B2 R2R_20k_0.B3 0.722031f
C77 D4 D3 0.115521f
C78 D5 V_REF 2.31749f
C79 a_1074_n2638# a_1776_n2638# 2.26e-19
C80 R2R_20k_0.B2 R2R_20k_0.B1 0.7282f
C81 a_n798_n2638# a_372_n2638# 1.94e-20
C82 a_2478_n2638# a_2244_n838# 0.401311f
C83 a_3648_n838# D6 0.001306f
C84 D1 a_138_n838# 0.001529f
C85 D3 V_REF 2.31853f
C86 a_2244_n838# R2R_20k_0.B5 2.11e-20
C87 R2R_20k_0.B7 a_3648_n838# 1.19e-20
C88 D3 a_1542_n838# 0.001537f
C89 a_n564_n838# a_n798_n2638# 0.006309f
C90 R2R_20k_0.B6 V_REF 5.80222f
C91 D4 R2R_20k_0.B5 1.99e-19
C92 R2R_20k_0.B3 a_1776_n2638# 0.002521f
C93 R2R_20k_0.B7 V_out 0.772359f
C94 R2R_20k_0.B2 a_840_n838# 0.422662f
C95 a_372_n2638# a_n330_n2638# 3.04e-19
C96 a_1074_n2638# a_138_n838# 0.299348f
C97 a_3648_n838# a_2946_n838# 0.129383f
C98 a_2478_n2638# a_1542_n838# 0.296855f
C99 D1 D2 0.115519f
C100 D5 R2R_20k_0.B6 1.99e-19
C101 D7 V_REF 2.30714f
C102 R2R_20k_0.B5 V_REF 5.80222f
C103 a_n564_n838# a_n330_n2638# 0.400342f
C104 a_372_n2638# a_1776_n2638# 1.25e-20
C105 a_2946_n838# V_out 2.92e-20
C106 a_3180_n2638# a_2946_n838# 0.400577f
C107 R2R_20k_0.B2 V_REF 5.80222f
C108 R2R_20k_0.B2 R2R_20k_0.B0 8.1e-21
C109 R2R_20k_0.B2 a_1542_n838# 0.299129f
C110 D0 D2 3.9e-20
C111 R2R_20k_0.B7 D6 1.99e-19
C112 a_2244_n838# a_1776_n2638# 5.96e-21
C113 V_out R2R_20k_0.B4 5.68e-21
C114 a_840_n838# a_1776_n2638# 0.299386f
C115 D5 R2R_20k_0.B5 4.25458f
C116 a_3882_n2638# a_3648_n838# 0.40049f
C117 a_3648_n838# R2R_20k_0.B3 1.94e-21
C118 m4_n961_5637# D1 0.001155f
C119 R2R_20k_0.B1 a_138_n838# 0.447872f
C120 R2R_20k_0.B0 a_n330_n2638# 0.002521f
C121 a_372_n2638# a_138_n838# 0.401867f
C122 R2R_20k_0.B3 D2 1.99e-19
C123 m4_n961_5637# D0 0.008711f
C124 a_n564_n838# a_138_n838# 0.126023f
C125 D7 R2R_20k_0.B6 0.016236f
C126 R2R_20k_0.B5 R2R_20k_0.B6 0.709935f
C127 a_1542_n838# a_1776_n2638# 0.40112f
C128 a_840_n838# a_138_n838# 0.126468f
C129 R2R_20k_0.B2 D3 0.016236f
C130 R2R_20k_0.B1 D2 0.016236f
C131 D1 D0 0.116931f
C132 a_2946_n838# R2R_20k_0.B4 0.298874f
C133 R2R_20k_0.B0 a_138_n838# 0.29912f
C134 a_840_n838# D2 0.00168f
C135 a_3180_n2638# a_2244_n838# 0.297634f
C136 a_3882_n2638# a_2946_n838# 0.297431f
C137 a_2946_n838# R2R_20k_0.B3 2.6e-20
C138 V_out V_COM 1.38016f
C139 D7 V_COM 2.31677f
C140 D6 V_COM 2.180716f
C141 D5 V_COM 2.191726f
C142 D4 V_COM 2.191964f
C143 D3 V_COM 2.191819f
C144 D2 V_COM 2.191829f
C145 D1 V_COM 2.181076f
C146 D0 V_COM 2.343576f
C147 V_REF V_COM 78.41346f
C148 m4_n961_5637# V_COM 0.13949f $ **FLOATING
C149 a_4584_n2638# V_COM 0.918344f
C150 a_3882_n2638# V_COM 0.570951f
C151 a_3648_n838# V_COM 1.32139f
C152 a_3180_n2638# V_COM 0.571287f
C153 a_2946_n838# V_COM 1.20795f
C154 a_2478_n2638# V_COM 0.570697f
C155 a_2244_n838# V_COM 1.20818f
C156 a_1776_n2638# V_COM 0.573523f
C157 a_1542_n838# V_COM 1.20705f
C158 a_1074_n2638# V_COM 0.574167f
C159 a_840_n838# V_COM 1.20846f
C160 a_372_n2638# V_COM 0.579198f
C161 a_138_n838# V_COM 1.20996f
C162 a_n330_n2638# V_COM 0.573636f
C163 a_n564_n838# V_COM 1.61447f
C164 a_n798_n2638# V_COM 0.924823f
C165 R2R_20k_0.B7 V_COM 7.636687f
C166 R2R_20k_0.B6 V_COM 5.682888f
C167 R2R_20k_0.B5 V_COM 5.953592f
C168 R2R_20k_0.B4 V_COM 5.750403f
C169 R2R_20k_0.B3 V_COM 6.037802f
C170 R2R_20k_0.B2 V_COM 5.7629f
C171 R2R_20k_0.B1 V_COM 6.096395f
C172 R2R_20k_0.B0 V_COM 6.913474f
C173 R2R_20k_0.B3.t5 V_COM 0.17916f
C174 R2R_20k_0.B3.t4 V_COM 0.17916f
C175 R2R_20k_0.B3.n0 V_COM 1.06496f
C176 R2R_20k_0.B3.t1 V_COM 0.078382f
C177 R2R_20k_0.B3.t2 V_COM 0.078382f
C178 R2R_20k_0.B3.n1 V_COM 0.178338f
C179 R2R_20k_0.B3.n2 V_COM 2.38605f
C180 R2R_20k_0.B3.t6 V_COM 1.31972f
C181 R2R_20k_0.B3.t3 V_COM 0.285838f
C182 R2R_20k_0.B3.n3 V_COM 2.53828f
C183 R2R_20k_0.B3.n4 V_COM 0.407859f
C184 R2R_20k_0.B3.t0 V_COM 0.083552f
C185 R2R_20k_0.B3.n5 V_COM 0.807666f
C186 D3.t4 V_COM 0.856565f
C187 D3.n0 V_COM 0.432352f
C188 D3.t1 V_COM 0.856565f
C189 D3.t0 V_COM 0.393621f
C190 D3.t3 V_COM 0.393621f
C191 D3.t2 V_COM 0.393621f
C192 D3.t5 V_COM 0.856565f
C193 D3.n1 V_COM 0.426051f
C194 D3.n2 V_COM 0.112805f
C195 D3.n3 V_COM 0.116115f
C196 D3.n4 V_COM 0.112805f
C197 D3.n5 V_COM 0.438773f
C198 D3.n6 V_COM 0.503232f
C199 D6.t2 V_COM 0.84393f
C200 D6.n0 V_COM 0.426566f
C201 D6.t1 V_COM 0.84393f
C202 D6.t3 V_COM 0.387815f
C203 D6.t5 V_COM 0.387815f
C204 D6.t4 V_COM 0.387815f
C205 D6.t0 V_COM 0.84393f
C206 D6.n1 V_COM 0.419766f
C207 D6.n2 V_COM 0.111141f
C208 D6.n3 V_COM 0.114402f
C209 D6.n4 V_COM 0.111141f
C210 D6.n5 V_COM 0.431273f
C211 D6.n6 V_COM 0.494011f
C212 R2R_20k_0.B2.t3 V_COM 1.32117f
C213 R2R_20k_0.B2.t2 V_COM 0.286153f
C214 R2R_20k_0.B2.n0 V_COM 2.54165f
C215 R2R_20k_0.B2.t4 V_COM 0.179357f
C216 R2R_20k_0.B2.t5 V_COM 0.179357f
C217 R2R_20k_0.B2.n1 V_COM 1.06613f
C218 R2R_20k_0.B2.t0 V_COM 0.078469f
C219 R2R_20k_0.B2.t1 V_COM 0.078469f
C220 R2R_20k_0.B2.n2 V_COM 0.178535f
C221 R2R_20k_0.B2.n3 V_COM 2.3835f
C222 R2R_20k_0.B2.n4 V_COM 0.698282f
C223 R2R_20k_0.B2.t6 V_COM 0.083546f
C224 R2R_20k_0.B2.n5 V_COM 0.800663f
C225 D2.t3 V_COM 0.856565f
C226 D2.n0 V_COM 0.432352f
C227 D2.t4 V_COM 0.856565f
C228 D2.t1 V_COM 0.393621f
C229 D2.t5 V_COM 0.393621f
C230 D2.t2 V_COM 0.393621f
C231 D2.t0 V_COM 0.856565f
C232 D2.n1 V_COM 0.426051f
C233 D2.n2 V_COM 0.112805f
C234 D2.n3 V_COM 0.116115f
C235 D2.n4 V_COM 0.112805f
C236 D2.n5 V_COM 0.438773f
C237 D2.n6 V_COM 0.503232f
C238 R2R_20k_0.B4.t6 V_COM 1.3247f
C239 R2R_20k_0.B4.t1 V_COM 0.286917f
C240 R2R_20k_0.B4.n0 V_COM 2.54868f
C241 R2R_20k_0.B4.t5 V_COM 0.179836f
C242 R2R_20k_0.B4.t4 V_COM 0.179836f
C243 R2R_20k_0.B4.n1 V_COM 1.06898f
C244 R2R_20k_0.B4.t2 V_COM 0.078678f
C245 R2R_20k_0.B4.t3 V_COM 0.078678f
C246 R2R_20k_0.B4.n2 V_COM 0.179012f
C247 R2R_20k_0.B4.n3 V_COM 2.38987f
C248 R2R_20k_0.B4.n4 V_COM 0.661136f
C249 R2R_20k_0.B4.t0 V_COM 0.083991f
C250 R2R_20k_0.B4.n5 V_COM 0.799643f
C251 D4.t1 V_COM 0.856478f
C252 D4.n0 V_COM 0.433443f
C253 D4.t0 V_COM 0.856478f
C254 D4.t4 V_COM 0.393581f
C255 D4.t3 V_COM 0.393581f
C256 D4.t2 V_COM 0.393581f
C257 D4.t5 V_COM 0.856478f
C258 D4.n1 V_COM 0.426008f
C259 D4.n2 V_COM 0.112793f
C260 D4.n3 V_COM 0.116103f
C261 D4.n4 V_COM 0.112793f
C262 D4.n5 V_COM 0.437679f
C263 D4.n6 V_COM 0.503661f
C264 R2R_20k_0.B6.t5 V_COM 0.083815f
C265 R2R_20k_0.B6.t2 V_COM 1.32161f
C266 R2R_20k_0.B6.t3 V_COM 0.286249f
C267 R2R_20k_0.B6.n0 V_COM 2.54258f
C268 R2R_20k_0.B6.t6 V_COM 0.179417f
C269 R2R_20k_0.B6.t4 V_COM 0.179417f
C270 R2R_20k_0.B6.n1 V_COM 1.06649f
C271 R2R_20k_0.B6.t0 V_COM 0.078495f
C272 R2R_20k_0.B6.t1 V_COM 0.078495f
C273 R2R_20k_0.B6.n2 V_COM 0.178595f
C274 R2R_20k_0.B6.n3 V_COM 2.3843f
C275 R2R_20k_0.B6.n4 V_COM 0.606654f
C276 R2R_20k_0.B6.n5 V_COM 0.772834f
C277 R2R_20k_0.B7.t0 V_COM 0.077069f
C278 R2R_20k_0.B7.t5 V_COM 1.21524f
C279 R2R_20k_0.B7.t3 V_COM 0.26321f
C280 R2R_20k_0.B7.n0 V_COM 2.33301f
C281 R2R_20k_0.B7.t6 V_COM 0.164977f
C282 R2R_20k_0.B7.t4 V_COM 0.164977f
C283 R2R_20k_0.B7.n1 V_COM 0.980655f
C284 R2R_20k_0.B7.t1 V_COM 0.072177f
C285 R2R_20k_0.B7.t2 V_COM 0.072177f
C286 R2R_20k_0.B7.n2 V_COM 0.16422f
C287 R2R_20k_0.B7.n3 V_COM 2.1924f
C288 R2R_20k_0.B7.n4 V_COM 0.458822f
C289 R2R_20k_0.B7.n5 V_COM 0.693191f
C290 D7.t2 V_COM 0.843672f
C291 D7.n0 V_COM 0.425357f
C292 D7.t3 V_COM 0.843672f
C293 D7.t0 V_COM 0.387696f
C294 D7.t5 V_COM 0.387696f
C295 D7.t1 V_COM 0.387696f
C296 D7.t4 V_COM 0.843672f
C297 D7.n1 V_COM 0.419638f
C298 D7.n2 V_COM 0.111107f
C299 D7.n3 V_COM 0.114368f
C300 D7.n4 V_COM 0.111107f
C301 D7.n5 V_COM 0.432559f
C302 D7.n6 V_COM 0.495198f
C303 R2R_20k_0.B5.t6 V_COM 0.084374f
C304 R2R_20k_0.B5.t5 V_COM 0.180533f
C305 R2R_20k_0.B5.t3 V_COM 0.180533f
C306 R2R_20k_0.B5.n0 V_COM 1.07313f
C307 R2R_20k_0.B5.t2 V_COM 0.078983f
C308 R2R_20k_0.B5.t0 V_COM 0.078983f
C309 R2R_20k_0.B5.n1 V_COM 0.179706f
C310 R2R_20k_0.B5.n2 V_COM 2.40421f
C311 R2R_20k_0.B5.t4 V_COM 1.32983f
C312 R2R_20k_0.B5.t1 V_COM 0.288029f
C313 R2R_20k_0.B5.n3 V_COM 2.55774f
C314 R2R_20k_0.B5.n4 V_COM 0.411513f
C315 R2R_20k_0.B5.n5 V_COM 0.787461f
C316 D5.t0 V_COM 0.856652f
C317 D5.n0 V_COM 0.433183f
C318 D5.t1 V_COM 0.856652f
C319 D5.t4 V_COM 0.393661f
C320 D5.t2 V_COM 0.393661f
C321 D5.t5 V_COM 0.393661f
C322 D5.t3 V_COM 0.856652f
C323 D5.n1 V_COM 0.426094f
C324 D5.n2 V_COM 0.112816f
C325 D5.n3 V_COM 0.116127f
C326 D5.n4 V_COM 0.112816f
C327 D5.n5 V_COM 0.437897f
C328 D5.n6 V_COM 0.502852f
C329 R2R_20k_0.B0.t4 V_COM 0.179317f
C330 R2R_20k_0.B0.t6 V_COM 0.179317f
C331 R2R_20k_0.B0.n0 V_COM 1.0659f
C332 R2R_20k_0.B0.t1 V_COM 0.078451f
C333 R2R_20k_0.B0.t3 V_COM 0.078451f
C334 R2R_20k_0.B0.n1 V_COM 0.178495f
C335 R2R_20k_0.B0.n2 V_COM 2.38801f
C336 R2R_20k_0.B0.t5 V_COM 1.32088f
C337 R2R_20k_0.B0.t2 V_COM 0.286089f
C338 R2R_20k_0.B0.n3 V_COM 2.54051f
C339 R2R_20k_0.B0.n4 V_COM 0.40874f
C340 R2R_20k_0.B0.t0 V_COM 0.083637f
C341 R2R_20k_0.B0.n5 V_COM 0.837257f
C342 D0.t3 V_COM 0.876221f
C343 D0.n0 V_COM 0.447868f
C344 D0.t1 V_COM 0.876221f
C345 D0.t4 V_COM 0.402654f
C346 D0.t5 V_COM 0.402654f
C347 D0.t2 V_COM 0.402654f
C348 D0.t0 V_COM 0.876221f
C349 D0.n1 V_COM 0.435828f
C350 D0.n2 V_COM 0.115394f
C351 D0.n3 V_COM 0.11878f
C352 D0.n4 V_COM 0.115394f
C353 D0.n5 V_COM 0.444331f
C354 D0.n6 V_COM 0.531906f
C355 V_REF.t15 V_COM 0.415634f
C356 V_REF.t23 V_COM 0.084805f
C357 V_REF.t7 V_COM 0.084805f
C358 V_REF.n0 V_COM 0.279386f
C359 V_REF.n1 V_COM 0.477983f
C360 V_REF.n2 V_COM 0.232984f
C361 V_REF.n3 V_COM 0.239084f
C362 V_REF.t38 V_COM 1.98745f
C363 V_REF.n4 V_COM -5.94e-19
C364 V_REF.n5 V_COM 0.223568f
C365 V_REF.t39 V_COM 0.084805f
C366 V_REF.t43 V_COM 0.084805f
C367 V_REF.n6 V_COM 0.279386f
C368 V_REF.t25 V_COM 0.415748f
C369 V_REF.t5 V_COM 0.084805f
C370 V_REF.t13 V_COM 0.084805f
C371 V_REF.n7 V_COM 0.279386f
C372 V_REF.n8 V_COM 0.478019f
C373 V_REF.n9 V_COM 0.223568f
C374 V_REF.t4 V_COM 1.98745f
C375 V_REF.t24 V_COM 1.98745f
C376 V_REF.n10 V_COM 0.223568f
C377 V_REF.t2 V_COM 1.98745f
C378 V_REF.t34 V_COM 1.98745f
C379 V_REF.n11 V_COM 0.223568f
C380 V_REF.t3 V_COM 0.084805f
C381 V_REF.t1 V_COM 0.084805f
C382 V_REF.n12 V_COM 0.279386f
C383 V_REF.t45 V_COM 0.415748f
C384 V_REF.t11 V_COM 0.084805f
C385 V_REF.t37 V_COM 0.084805f
C386 V_REF.n13 V_COM 0.279386f
C387 V_REF.n14 V_COM 0.478019f
C388 V_REF.n15 V_COM 0.223568f
C389 V_REF.t10 V_COM 1.98745f
C390 V_REF.t44 V_COM 1.98745f
C391 V_REF.n16 V_COM 0.223568f
C392 V_REF.t20 V_COM 1.98745f
C393 V_REF.t18 V_COM 1.98745f
C394 V_REF.n17 V_COM 0.223568f
C395 V_REF.t21 V_COM 0.084805f
C396 V_REF.t9 V_COM 0.084805f
C397 V_REF.n18 V_COM 0.279386f
C398 V_REF.t27 V_COM 0.415748f
C399 V_REF.t17 V_COM 0.084805f
C400 V_REF.t33 V_COM 0.084805f
C401 V_REF.n19 V_COM 0.279386f
C402 V_REF.n20 V_COM 0.478019f
C403 V_REF.n21 V_COM 0.223568f
C404 V_REF.t16 V_COM 1.98745f
C405 V_REF.t26 V_COM 1.98745f
C406 V_REF.t29 V_COM 0.084805f
C407 V_REF.t47 V_COM 0.084805f
C408 V_REF.n22 V_COM 0.28057f
C409 V_REF.t31 V_COM 0.415748f
C410 V_REF.n23 V_COM 0.53035f
C411 V_REF.n24 V_COM 0.88405f
C412 V_REF.n25 V_COM 0.248138f
C413 V_REF.t28 V_COM 2.63406f
C414 V_REF.t30 V_COM 1.98745f
C415 V_REF.t46 V_COM 1.0754f
C416 V_REF.n26 V_COM 0.202351f
C417 V_REF.n27 V_COM 0.229244f
C418 V_REF.n28 V_COM 0.001049f
C419 V_REF.t32 V_COM 1.0754f
C420 V_REF.n29 V_COM 0.041161f
C421 V_REF.n30 V_COM 0.140407f
C422 V_REF.n31 V_COM 0.53035f
C423 V_REF.n32 V_COM 0.478019f
C424 V_REF.t19 V_COM 0.415748f
C425 V_REF.n33 V_COM 0.53035f
C426 V_REF.n34 V_COM 0.140407f
C427 V_REF.n35 V_COM 0.041161f
C428 V_REF.t8 V_COM 1.0754f
C429 V_REF.n36 V_COM 0.001049f
C430 V_REF.n37 V_COM 0.223568f
C431 V_REF.n38 V_COM 0.001049f
C432 V_REF.t36 V_COM 1.0754f
C433 V_REF.n39 V_COM 0.041161f
C434 V_REF.n40 V_COM 0.140407f
C435 V_REF.n41 V_COM 0.53035f
C436 V_REF.n42 V_COM 0.478019f
C437 V_REF.t35 V_COM 0.415748f
C438 V_REF.n43 V_COM 0.53035f
C439 V_REF.n44 V_COM 0.140407f
C440 V_REF.n45 V_COM 0.041161f
C441 V_REF.t0 V_COM 1.0754f
C442 V_REF.n46 V_COM 0.001049f
C443 V_REF.n47 V_COM 0.223568f
C444 V_REF.n48 V_COM 0.223568f
C445 V_REF.n49 V_COM 0.001049f
C446 V_REF.t12 V_COM 1.0754f
C447 V_REF.n50 V_COM 0.041161f
C448 V_REF.n51 V_COM 0.140407f
C449 V_REF.n52 V_COM 0.53035f
C450 V_REF.n53 V_COM 0.478019f
C451 V_REF.t41 V_COM 0.415748f
C452 V_REF.n54 V_COM 0.073474f
C453 V_REF.n55 V_COM 0.51061f
C454 V_REF.n56 V_COM 0.140407f
C455 V_REF.n57 V_COM 0.039638f
C456 V_REF.t42 V_COM 1.0754f
C457 V_REF.t40 V_COM 1.98092f
C458 V_REF.t22 V_COM 1.98108f
C459 V_REF.t14 V_COM 2.63406f
C460 V_REF.t6 V_COM 1.0754f
C461 V_REF.n58 V_COM 0.200405f
C462 V_REF.n59 V_COM 0.246495f
C463 V_REF.n60 V_COM 0.140935f
C464 V_REF.n61 V_COM 0.531655f
C465 R2R_20k_0.B1.t1 V_COM 0.176173f
C466 R2R_20k_0.B1.t2 V_COM 0.176173f
C467 R2R_20k_0.B1.n0 V_COM 1.04721f
C468 R2R_20k_0.B1.t5 V_COM 0.077076f
C469 R2R_20k_0.B1.t0 V_COM 0.077076f
C470 R2R_20k_0.B1.n1 V_COM 0.175365f
C471 R2R_20k_0.B1.n2 V_COM 2.34628f
C472 R2R_20k_0.B1.t3 V_COM 1.29772f
C473 R2R_20k_0.B1.t4 V_COM 0.281073f
C474 R2R_20k_0.B1.n3 V_COM 2.49581f
C475 R2R_20k_0.B1.n4 V_COM 0.401593f
C476 R2R_20k_0.B1.t6 V_COM 0.082044f
C477 R2R_20k_0.B1.n5 V_COM 0.822102f
C478 D1.t0 V_COM 0.843844f
C479 D1.n0 V_COM 0.425099f
C480 D1.t3 V_COM 0.843844f
C481 D1.t4 V_COM 0.387775f
C482 D1.t5 V_COM 0.387775f
C483 D1.t1 V_COM 0.387775f
C484 D1.t2 V_COM 0.843844f
C485 D1.n1 V_COM 0.419724f
C486 D1.n2 V_COM 0.11113f
C487 D1.n3 V_COM 0.114391f
C488 D1.n4 V_COM 0.11113f
C489 D1.n5 V_COM 0.432786f
C490 D1.n6 V_COM 0.494387f
.ends

