** sch_path: /home/ttuser/tinytapeout/TT_Project/xschem/sar_adc_analog.sch
.subckt sar_adc_analog SH V_in comp_out ibias D0 VDDA D1 D2 D3 VSSA D4 V_REF D5 D6 D7 v_sh_out dac_out
*.PININFO D0:I comp_out:O D1:I D2:I D3:I D4:I D5:I D6:I D7:I V_REF:I SH:I V_in:I VDDA:I VSSA:I ibias:I dac_out:O v_sh_out:O
x1 dac_out D7 D0 D1 D6 D2 D5 D3 D4 V_REF VSSA r2r_dac
x2 VDDA ibias v_sh_out dac_out comp_out VSSA comparator
x3 VDDA SH v_sh_out V_in VSSA sample_hold
.ends

* expanding   symbol:  r2r_dac.sym # of pins=11
** sym_path: /home/ttuser/tinytapeout/TT_Project/xschem/r2r_dac.sym
** sch_path: /home/ttuser/tinytapeout/TT_Project/xschem/r2r_dac.sch
.subckt r2r_dac V_out D7 D0 D1 D6 D2 D5 D3 D4 V_REF V_COM
*.PININFO D0:I V_out:O V_REF:B V_COM:B D1:I D2:I D3:I D7:I D6:I D5:I D4:I
x1 net2 net1 net3 net4 net8 net5 net7 net6 V_COM V_out R2R_20k
x2 V_REF D0 net1 V_COM dac_switch
x3 V_REF D1 net2 V_COM dac_switch
x4 V_REF D2 net3 V_COM dac_switch
x5 V_REF D3 net4 V_COM dac_switch
x6 V_REF D7 net8 V_COM dac_switch
x7 V_REF D6 net7 V_COM dac_switch
x8 V_REF D5 net6 V_COM dac_switch
x9 V_REF D4 net5 V_COM dac_switch
.ends
meas tran b1_logic FIND v(v_b1) AT=10n THRESHOLD=0.5

* expanding   symbol:  comparator.sym # of pins=6
** sym_path: /home/ttuser/tinytapeout/TT_Project/xschem/comparator.sym
** sch_path: /home/ttuser/tinytapeout/TT_Project/xschem/comparator.sch
.subckt comparator vdda ibias inp inn outp vssa
*.PININFO ibias:I inn:I inp:I outp:O vdda:I vssa:I
XM1[1] vsp ibias vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=8 m=1
XM1[2] vsp ibias vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=8 m=1
XM2 ibias ibias vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=8 m=1
XM3[1] vgsn inn vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM3[2] vgsn inn vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM3[3] vgsn inn vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM3[4] vgsn inn vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM4[1] vout1 inp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM4[2] vout1 inp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM4[3] vout1 inp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM4[4] vout1 inp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=2 m=1
XM5[1] vout1 vgsn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=1 W=18 nf=2 m=1
XM5[2] vout1 vgsn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=1 W=18 nf=2 m=1
XM6[1] vgsn vgsn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=1 W=18 nf=2 m=1
XM6[2] vgsn vgsn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=1 W=18 nf=2 m=1
XM7 outp voutinv1 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM8 outp voutinv1 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM9 vout2 vout1 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=1 W=70 nf=4 m=1
XM10[1] vout2 ibias vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=8 m=1
XM10[2] vout2 ibias vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=50 nf=8 m=1
XM11 voutinv1 vout2 vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=1 m=1
XM12 voutinv1 vout2 vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XMDY3[1] vssa vgsn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=1 W=9 nf=2 m=1
XMDY3[2] vssa vgsn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=1 W=9 nf=2 m=1
XMDY1[1] vdda ibias vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=8 m=1
XMDY1[2] vdda ibias vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=20 nf=8 m=1
XMDY2[1] vsp vsp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=25 nf=1 m=1
XMDY2[2] vsp vsp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=25 nf=1 m=1
XMDY2[3] vsp vsp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=25 nf=1 m=1
XMDY2[4] vsp vsp vsp vdda sky130_fd_pr__pfet_g5v0d10v5 L=1 W=25 nf=1 m=1
.ends


* expanding   symbol:  sample_hold.sym # of pins=5
** sym_path: /home/ttuser/tinytapeout/TT_Project/xschem/sample_hold.sym
** sch_path: /home/ttuser/tinytapeout/TT_Project/xschem/sample_hold.sch
.subckt sample_hold vdda sample vout vin vssa
*.PININFO vout:O vdda:I vssa:I vin:I sample:I
XM5 vout sample vin vssa sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 nf=1 m=1
XM6 vout sample_n vin vdda sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=30 nf=3 m=1
XM3 sample_n sample vssa vssa sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM4 sample_n sample vdda vdda sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 nf=3 m=1
XC1 vout vssa sky130_fd_pr__cap_mim_m3_1 W=17 L=30 m=1
.ends


* expanding   symbol:  R2R_20k.sym # of pins=10
** sym_path: /home/ttuser/tinytapeout/TT_Project/xschem/R2R_20k.sym
** sch_path: /home/ttuser/tinytapeout/TT_Project/xschem/R2R_20k.sch
.subckt R2R_20k B1 B0 B2 B3 B7 B4 B6 B5 COM OUT
*.PININFO COM:B B0:B B1:B OUT:B B2:B B3:B B4:B B5:B B6:B B7:B
XR1 net1 H COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR2 B3 net1 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR3 net2 net13 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR4 B4 net2 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR5 net3 net14 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR6 B5 net3 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR7 net4 net15 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR8 B6 net4 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR9 net5 net9 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR10 COM net5 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR11 net6 net9 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR12 B0 net6 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR13 net7 net10 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR14 B1 net7 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR15 net8 net11 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR16 B2 net8 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR18 net10 net9 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR19 net11 net10 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR20 net13 H COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR21 net14 net13 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR22 net15 net14 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR17 net12 OUT COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR23 B7 net12 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR24 OUT net15 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR25 H net11 COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR26 COM COM COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
XR27 COM COM COM sky130_fd_pr__res_xhigh_po_0p69 L=7 mult=1 m=1
.ends


* expanding   symbol:  dac_switch.sym # of pins=4
** sym_path: /home/ttuser/tinytapeout/TT_Project/xschem/dac_switch.sym
** sch_path: /home/ttuser/tinytapeout/TT_Project/xschem/dac_switch.sch
.subckt dac_switch Vref Dx Outx Vcom
*.PININFO Dx:I Outx:O Vref:B Vcom:B
XM1 Outx Dx Vref Vref sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=48 nf=3 m=1
XM2 Outx Dx Vcom Vcom sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=21 nf=3 m=1
.ends

.end
