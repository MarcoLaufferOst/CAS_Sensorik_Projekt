magic
tech sky130A
magscale 1 2
timestamp 1736061100
<< error_p >>
rect -1127 -691 -1097 691
rect -1061 -625 -1031 625
rect 1031 -625 1061 625
rect 1097 -691 1127 691
<< nwell >>
rect -1097 -725 1097 725
<< mvpmos >>
rect -1003 -625 -803 625
rect -745 -625 -545 625
rect -487 -625 -287 625
rect -229 -625 -29 625
rect 29 -625 229 625
rect 287 -625 487 625
rect 545 -625 745 625
rect 803 -625 1003 625
<< mvpdiff >>
rect -1061 613 -1003 625
rect -1061 -613 -1049 613
rect -1015 -613 -1003 613
rect -1061 -625 -1003 -613
rect -803 613 -745 625
rect -803 -613 -791 613
rect -757 -613 -745 613
rect -803 -625 -745 -613
rect -545 613 -487 625
rect -545 -613 -533 613
rect -499 -613 -487 613
rect -545 -625 -487 -613
rect -287 613 -229 625
rect -287 -613 -275 613
rect -241 -613 -229 613
rect -287 -625 -229 -613
rect -29 613 29 625
rect -29 -613 -17 613
rect 17 -613 29 613
rect -29 -625 29 -613
rect 229 613 287 625
rect 229 -613 241 613
rect 275 -613 287 613
rect 229 -625 287 -613
rect 487 613 545 625
rect 487 -613 499 613
rect 533 -613 545 613
rect 487 -625 545 -613
rect 745 613 803 625
rect 745 -613 757 613
rect 791 -613 803 613
rect 745 -625 803 -613
rect 1003 613 1061 625
rect 1003 -613 1015 613
rect 1049 -613 1061 613
rect 1003 -625 1061 -613
<< mvpdiffc >>
rect -1049 -613 -1015 613
rect -791 -613 -757 613
rect -533 -613 -499 613
rect -275 -613 -241 613
rect -17 -613 17 613
rect 241 -613 275 613
rect 499 -613 533 613
rect 757 -613 791 613
rect 1015 -613 1049 613
<< poly >>
rect -1003 706 -803 722
rect -1003 672 -987 706
rect -819 672 -803 706
rect -1003 625 -803 672
rect -745 706 -545 722
rect -745 672 -729 706
rect -561 672 -545 706
rect -745 625 -545 672
rect -487 706 -287 722
rect -487 672 -471 706
rect -303 672 -287 706
rect -487 625 -287 672
rect -229 706 -29 722
rect -229 672 -213 706
rect -45 672 -29 706
rect -229 625 -29 672
rect 29 706 229 722
rect 29 672 45 706
rect 213 672 229 706
rect 29 625 229 672
rect 287 706 487 722
rect 287 672 303 706
rect 471 672 487 706
rect 287 625 487 672
rect 545 706 745 722
rect 545 672 561 706
rect 729 672 745 706
rect 545 625 745 672
rect 803 706 1003 722
rect 803 672 819 706
rect 987 672 1003 706
rect 803 625 1003 672
rect -1003 -672 -803 -625
rect -1003 -706 -987 -672
rect -819 -706 -803 -672
rect -1003 -722 -803 -706
rect -745 -672 -545 -625
rect -745 -706 -729 -672
rect -561 -706 -545 -672
rect -745 -722 -545 -706
rect -487 -672 -287 -625
rect -487 -706 -471 -672
rect -303 -706 -287 -672
rect -487 -722 -287 -706
rect -229 -672 -29 -625
rect -229 -706 -213 -672
rect -45 -706 -29 -672
rect -229 -722 -29 -706
rect 29 -672 229 -625
rect 29 -706 45 -672
rect 213 -706 229 -672
rect 29 -722 229 -706
rect 287 -672 487 -625
rect 287 -706 303 -672
rect 471 -706 487 -672
rect 287 -722 487 -706
rect 545 -672 745 -625
rect 545 -706 561 -672
rect 729 -706 745 -672
rect 545 -722 745 -706
rect 803 -672 1003 -625
rect 803 -706 819 -672
rect 987 -706 1003 -672
rect 803 -722 1003 -706
<< polycont >>
rect -987 672 -819 706
rect -729 672 -561 706
rect -471 672 -303 706
rect -213 672 -45 706
rect 45 672 213 706
rect 303 672 471 706
rect 561 672 729 706
rect 819 672 987 706
rect -987 -706 -819 -672
rect -729 -706 -561 -672
rect -471 -706 -303 -672
rect -213 -706 -45 -672
rect 45 -706 213 -672
rect 303 -706 471 -672
rect 561 -706 729 -672
rect 819 -706 987 -672
<< locali >>
rect -1003 672 -987 706
rect -819 672 -803 706
rect -745 672 -729 706
rect -561 672 -545 706
rect -487 672 -471 706
rect -303 672 -287 706
rect -229 672 -213 706
rect -45 672 -29 706
rect 29 672 45 706
rect 213 672 229 706
rect 287 672 303 706
rect 471 672 487 706
rect 545 672 561 706
rect 729 672 745 706
rect 803 672 819 706
rect 987 672 1003 706
rect -1049 613 -1015 629
rect -1049 -629 -1015 -613
rect -791 613 -757 629
rect -791 -629 -757 -613
rect -533 613 -499 629
rect -533 -629 -499 -613
rect -275 613 -241 629
rect -275 -629 -241 -613
rect -17 613 17 629
rect -17 -629 17 -613
rect 241 613 275 629
rect 241 -629 275 -613
rect 499 613 533 629
rect 499 -629 533 -613
rect 757 613 791 629
rect 757 -629 791 -613
rect 1015 613 1049 629
rect 1015 -629 1049 -613
rect -1003 -706 -987 -672
rect -819 -706 -803 -672
rect -745 -706 -729 -672
rect -561 -706 -545 -672
rect -487 -706 -471 -672
rect -303 -706 -287 -672
rect -229 -706 -213 -672
rect -45 -706 -29 -672
rect 29 -706 45 -672
rect 213 -706 229 -672
rect 287 -706 303 -672
rect 471 -706 487 -672
rect 545 -706 561 -672
rect 729 -706 745 -672
rect 803 -706 819 -672
rect 987 -706 1003 -672
<< viali >>
rect -987 672 -819 706
rect -729 672 -561 706
rect -471 672 -303 706
rect -213 672 -45 706
rect 45 672 213 706
rect 303 672 471 706
rect 561 672 729 706
rect 819 672 987 706
rect -1049 -613 -1015 613
rect -791 -613 -757 613
rect -533 -613 -499 613
rect -275 -613 -241 613
rect -17 -613 17 613
rect 241 -613 275 613
rect 499 -613 533 613
rect 757 -613 791 613
rect 1015 -613 1049 613
rect -987 -706 -819 -672
rect -729 -706 -561 -672
rect -471 -706 -303 -672
rect -213 -706 -45 -672
rect 45 -706 213 -672
rect 303 -706 471 -672
rect 561 -706 729 -672
rect 819 -706 987 -672
<< metal1 >>
rect -999 706 -807 712
rect -999 672 -987 706
rect -819 672 -807 706
rect -999 666 -807 672
rect -741 706 -549 712
rect -741 672 -729 706
rect -561 672 -549 706
rect -741 666 -549 672
rect -483 706 -291 712
rect -483 672 -471 706
rect -303 672 -291 706
rect -483 666 -291 672
rect -225 706 -33 712
rect -225 672 -213 706
rect -45 672 -33 706
rect -225 666 -33 672
rect 33 706 225 712
rect 33 672 45 706
rect 213 672 225 706
rect 33 666 225 672
rect 291 706 483 712
rect 291 672 303 706
rect 471 672 483 706
rect 291 666 483 672
rect 549 706 741 712
rect 549 672 561 706
rect 729 672 741 706
rect 549 666 741 672
rect 807 706 999 712
rect 807 672 819 706
rect 987 672 999 706
rect 807 666 999 672
rect -1055 613 -1009 625
rect -1055 -613 -1049 613
rect -1015 -613 -1009 613
rect -1055 -625 -1009 -613
rect -797 613 -751 625
rect -797 -613 -791 613
rect -757 -613 -751 613
rect -797 -625 -751 -613
rect -539 613 -493 625
rect -539 -613 -533 613
rect -499 -613 -493 613
rect -539 -625 -493 -613
rect -281 613 -235 625
rect -281 -613 -275 613
rect -241 -613 -235 613
rect -281 -625 -235 -613
rect -23 613 23 625
rect -23 -613 -17 613
rect 17 -613 23 613
rect -23 -625 23 -613
rect 235 613 281 625
rect 235 -613 241 613
rect 275 -613 281 613
rect 235 -625 281 -613
rect 493 613 539 625
rect 493 -613 499 613
rect 533 -613 539 613
rect 493 -625 539 -613
rect 751 613 797 625
rect 751 -613 757 613
rect 791 -613 797 613
rect 751 -625 797 -613
rect 1009 613 1055 625
rect 1009 -613 1015 613
rect 1049 -613 1055 613
rect 1009 -625 1055 -613
rect -999 -672 -807 -666
rect -999 -706 -987 -672
rect -819 -706 -807 -672
rect -999 -712 -807 -706
rect -741 -672 -549 -666
rect -741 -706 -729 -672
rect -561 -706 -549 -672
rect -741 -712 -549 -706
rect -483 -672 -291 -666
rect -483 -706 -471 -672
rect -303 -706 -291 -672
rect -483 -712 -291 -706
rect -225 -672 -33 -666
rect -225 -706 -213 -672
rect -45 -706 -33 -672
rect -225 -712 -33 -706
rect 33 -672 225 -666
rect 33 -706 45 -672
rect 213 -706 225 -672
rect 33 -712 225 -706
rect 291 -672 483 -666
rect 291 -706 303 -672
rect 471 -706 483 -672
rect 291 -712 483 -706
rect 549 -672 741 -666
rect 549 -706 561 -672
rect 729 -706 741 -672
rect 549 -712 741 -706
rect 807 -672 999 -666
rect 807 -706 819 -672
rect 987 -706 999 -672
rect 807 -712 999 -706
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6.25 l 1.0 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
