magic
tech sky130A
magscale 1 2
timestamp 1737184964
<< mvnmos >>
rect -1003 -1500 -803 1500
rect -745 -1500 -545 1500
rect -487 -1500 -287 1500
rect -229 -1500 -29 1500
rect 29 -1500 229 1500
rect 287 -1500 487 1500
rect 545 -1500 745 1500
rect 803 -1500 1003 1500
<< mvndiff >>
rect -1061 1488 -1003 1500
rect -1061 -1488 -1049 1488
rect -1015 -1488 -1003 1488
rect -1061 -1500 -1003 -1488
rect -803 1488 -745 1500
rect -803 -1488 -791 1488
rect -757 -1488 -745 1488
rect -803 -1500 -745 -1488
rect -545 1488 -487 1500
rect -545 -1488 -533 1488
rect -499 -1488 -487 1488
rect -545 -1500 -487 -1488
rect -287 1488 -229 1500
rect -287 -1488 -275 1488
rect -241 -1488 -229 1488
rect -287 -1500 -229 -1488
rect -29 1488 29 1500
rect -29 -1488 -17 1488
rect 17 -1488 29 1488
rect -29 -1500 29 -1488
rect 229 1488 287 1500
rect 229 -1488 241 1488
rect 275 -1488 287 1488
rect 229 -1500 287 -1488
rect 487 1488 545 1500
rect 487 -1488 499 1488
rect 533 -1488 545 1488
rect 487 -1500 545 -1488
rect 745 1488 803 1500
rect 745 -1488 757 1488
rect 791 -1488 803 1488
rect 745 -1500 803 -1488
rect 1003 1488 1061 1500
rect 1003 -1488 1015 1488
rect 1049 -1488 1061 1488
rect 1003 -1500 1061 -1488
<< mvndiffc >>
rect -1049 -1488 -1015 1488
rect -791 -1488 -757 1488
rect -533 -1488 -499 1488
rect -275 -1488 -241 1488
rect -17 -1488 17 1488
rect 241 -1488 275 1488
rect 499 -1488 533 1488
rect 757 -1488 791 1488
rect 1015 -1488 1049 1488
<< poly >>
rect -1003 1572 -803 1588
rect -1003 1538 -987 1572
rect -819 1538 -803 1572
rect -1003 1500 -803 1538
rect -745 1572 -545 1588
rect -745 1538 -729 1572
rect -561 1538 -545 1572
rect -745 1500 -545 1538
rect -487 1572 -287 1588
rect -487 1538 -471 1572
rect -303 1538 -287 1572
rect -487 1500 -287 1538
rect -229 1572 -29 1588
rect -229 1538 -213 1572
rect -45 1538 -29 1572
rect -229 1500 -29 1538
rect 29 1572 229 1588
rect 29 1538 45 1572
rect 213 1538 229 1572
rect 29 1500 229 1538
rect 287 1572 487 1588
rect 287 1538 303 1572
rect 471 1538 487 1572
rect 287 1500 487 1538
rect 545 1572 745 1588
rect 545 1538 561 1572
rect 729 1538 745 1572
rect 545 1500 745 1538
rect 803 1572 1003 1588
rect 803 1538 819 1572
rect 987 1538 1003 1572
rect 803 1500 1003 1538
rect -1003 -1538 -803 -1500
rect -1003 -1572 -987 -1538
rect -819 -1572 -803 -1538
rect -1003 -1588 -803 -1572
rect -745 -1538 -545 -1500
rect -745 -1572 -729 -1538
rect -561 -1572 -545 -1538
rect -745 -1588 -545 -1572
rect -487 -1538 -287 -1500
rect -487 -1572 -471 -1538
rect -303 -1572 -287 -1538
rect -487 -1588 -287 -1572
rect -229 -1538 -29 -1500
rect -229 -1572 -213 -1538
rect -45 -1572 -29 -1538
rect -229 -1588 -29 -1572
rect 29 -1538 229 -1500
rect 29 -1572 45 -1538
rect 213 -1572 229 -1538
rect 29 -1588 229 -1572
rect 287 -1538 487 -1500
rect 287 -1572 303 -1538
rect 471 -1572 487 -1538
rect 287 -1588 487 -1572
rect 545 -1538 745 -1500
rect 545 -1572 561 -1538
rect 729 -1572 745 -1538
rect 545 -1588 745 -1572
rect 803 -1538 1003 -1500
rect 803 -1572 819 -1538
rect 987 -1572 1003 -1538
rect 803 -1588 1003 -1572
<< polycont >>
rect -987 1538 -819 1572
rect -729 1538 -561 1572
rect -471 1538 -303 1572
rect -213 1538 -45 1572
rect 45 1538 213 1572
rect 303 1538 471 1572
rect 561 1538 729 1572
rect 819 1538 987 1572
rect -987 -1572 -819 -1538
rect -729 -1572 -561 -1538
rect -471 -1572 -303 -1538
rect -213 -1572 -45 -1538
rect 45 -1572 213 -1538
rect 303 -1572 471 -1538
rect 561 -1572 729 -1538
rect 819 -1572 987 -1538
<< locali >>
rect -1003 1538 -987 1572
rect -819 1538 -803 1572
rect -745 1538 -729 1572
rect -561 1538 -545 1572
rect -487 1538 -471 1572
rect -303 1538 -287 1572
rect -229 1538 -213 1572
rect -45 1538 -29 1572
rect 29 1538 45 1572
rect 213 1538 229 1572
rect 287 1538 303 1572
rect 471 1538 487 1572
rect 545 1538 561 1572
rect 729 1538 745 1572
rect 803 1538 819 1572
rect 987 1538 1003 1572
rect -1049 1488 -1015 1504
rect -1049 -1504 -1015 -1488
rect -791 1488 -757 1504
rect -791 -1504 -757 -1488
rect -533 1488 -499 1504
rect -533 -1504 -499 -1488
rect -275 1488 -241 1504
rect -275 -1504 -241 -1488
rect -17 1488 17 1504
rect -17 -1504 17 -1488
rect 241 1488 275 1504
rect 241 -1504 275 -1488
rect 499 1488 533 1504
rect 499 -1504 533 -1488
rect 757 1488 791 1504
rect 757 -1504 791 -1488
rect 1015 1488 1049 1504
rect 1015 -1504 1049 -1488
rect -1003 -1572 -987 -1538
rect -819 -1572 -803 -1538
rect -745 -1572 -729 -1538
rect -561 -1572 -545 -1538
rect -487 -1572 -471 -1538
rect -303 -1572 -287 -1538
rect -229 -1572 -213 -1538
rect -45 -1572 -29 -1538
rect 29 -1572 45 -1538
rect 213 -1572 229 -1538
rect 287 -1572 303 -1538
rect 471 -1572 487 -1538
rect 545 -1572 561 -1538
rect 729 -1572 745 -1538
rect 803 -1572 819 -1538
rect 987 -1572 1003 -1538
<< viali >>
rect -987 1538 -819 1572
rect -729 1538 -561 1572
rect -471 1538 -303 1572
rect -213 1538 -45 1572
rect 45 1538 213 1572
rect 303 1538 471 1572
rect 561 1538 729 1572
rect 819 1538 987 1572
rect -1049 -1488 -1015 1488
rect -791 -1488 -757 1488
rect -533 -1488 -499 1488
rect -275 -1488 -241 1488
rect -17 -1488 17 1488
rect 241 -1488 275 1488
rect 499 -1488 533 1488
rect 757 -1488 791 1488
rect 1015 -1488 1049 1488
rect -987 -1572 -819 -1538
rect -729 -1572 -561 -1538
rect -471 -1572 -303 -1538
rect -213 -1572 -45 -1538
rect 45 -1572 213 -1538
rect 303 -1572 471 -1538
rect 561 -1572 729 -1538
rect 819 -1572 987 -1538
<< metal1 >>
rect -999 1572 -807 1578
rect -999 1538 -987 1572
rect -819 1538 -807 1572
rect -999 1532 -807 1538
rect -741 1572 -549 1578
rect -741 1538 -729 1572
rect -561 1538 -549 1572
rect -741 1532 -549 1538
rect -483 1572 -291 1578
rect -483 1538 -471 1572
rect -303 1538 -291 1572
rect -483 1532 -291 1538
rect -225 1572 -33 1578
rect -225 1538 -213 1572
rect -45 1538 -33 1572
rect -225 1532 -33 1538
rect 33 1572 225 1578
rect 33 1538 45 1572
rect 213 1538 225 1572
rect 33 1532 225 1538
rect 291 1572 483 1578
rect 291 1538 303 1572
rect 471 1538 483 1572
rect 291 1532 483 1538
rect 549 1572 741 1578
rect 549 1538 561 1572
rect 729 1538 741 1572
rect 549 1532 741 1538
rect 807 1572 999 1578
rect 807 1538 819 1572
rect 987 1538 999 1572
rect 807 1532 999 1538
rect -1055 1488 -1009 1500
rect -1055 -1488 -1049 1488
rect -1015 -1488 -1009 1488
rect -1055 -1500 -1009 -1488
rect -797 1488 -751 1500
rect -797 -1488 -791 1488
rect -757 -1488 -751 1488
rect -797 -1500 -751 -1488
rect -539 1488 -493 1500
rect -539 -1488 -533 1488
rect -499 -1488 -493 1488
rect -539 -1500 -493 -1488
rect -281 1488 -235 1500
rect -281 -1488 -275 1488
rect -241 -1488 -235 1488
rect -281 -1500 -235 -1488
rect -23 1488 23 1500
rect -23 -1488 -17 1488
rect 17 -1488 23 1488
rect -23 -1500 23 -1488
rect 235 1488 281 1500
rect 235 -1488 241 1488
rect 275 -1488 281 1488
rect 235 -1500 281 -1488
rect 493 1488 539 1500
rect 493 -1488 499 1488
rect 533 -1488 539 1488
rect 493 -1500 539 -1488
rect 751 1488 797 1500
rect 751 -1488 757 1488
rect 791 -1488 797 1488
rect 751 -1500 797 -1488
rect 1009 1488 1055 1500
rect 1009 -1488 1015 1488
rect 1049 -1488 1055 1488
rect 1009 -1500 1055 -1488
rect -999 -1538 -807 -1532
rect -999 -1572 -987 -1538
rect -819 -1572 -807 -1538
rect -999 -1578 -807 -1572
rect -741 -1538 -549 -1532
rect -741 -1572 -729 -1538
rect -561 -1572 -549 -1538
rect -741 -1578 -549 -1572
rect -483 -1538 -291 -1532
rect -483 -1572 -471 -1538
rect -303 -1572 -291 -1538
rect -483 -1578 -291 -1572
rect -225 -1538 -33 -1532
rect -225 -1572 -213 -1538
rect -45 -1572 -33 -1538
rect -225 -1578 -33 -1572
rect 33 -1538 225 -1532
rect 33 -1572 45 -1538
rect 213 -1572 225 -1538
rect 33 -1578 225 -1572
rect 291 -1538 483 -1532
rect 291 -1572 303 -1538
rect 471 -1572 483 -1538
rect 291 -1578 483 -1572
rect 549 -1538 741 -1532
rect 549 -1572 561 -1538
rect 729 -1572 741 -1538
rect 549 -1578 741 -1572
rect 807 -1538 999 -1532
rect 807 -1572 819 -1538
rect 987 -1572 999 -1538
rect 807 -1578 999 -1572
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 15 l 1 m 1 nf 8 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
