magic
tech sky130A
magscale 1 2
timestamp 1736113453
<< pwell >>
rect -3277 -1282 3277 1282
<< psubdiff >>
rect -3241 1212 3241 1246
rect -3241 1150 -3207 1212
rect 3207 1150 3241 1212
rect -3241 -1212 -3207 -1150
rect 3207 -1212 3241 -1150
rect -3241 -1246 -3145 -1212
rect 3145 -1246 3241 -1212
<< psubdiffcont >>
rect -3241 -1150 -3207 1150
rect 3207 -1150 3241 1150
rect -3145 -1246 3145 -1212
<< xpolycontact >>
rect -3111 684 -2973 1116
rect -3111 -1116 -2973 -684
rect -2877 684 -2739 1116
rect -2877 -1116 -2739 -684
rect -2643 684 -2505 1116
rect -2643 -1116 -2505 -684
rect -2409 684 -2271 1116
rect -2409 -1116 -2271 -684
rect -2175 684 -2037 1116
rect -2175 -1116 -2037 -684
rect -1941 684 -1803 1116
rect -1941 -1116 -1803 -684
rect -1707 684 -1569 1116
rect -1707 -1116 -1569 -684
rect -1473 684 -1335 1116
rect -1473 -1116 -1335 -684
rect -1239 684 -1101 1116
rect -1239 -1116 -1101 -684
rect -1005 684 -867 1116
rect -1005 -1116 -867 -684
rect -771 684 -633 1116
rect -771 -1116 -633 -684
rect -537 684 -399 1116
rect -537 -1116 -399 -684
rect -303 684 -165 1116
rect -303 -1116 -165 -684
rect -69 684 69 1116
rect -69 -1116 69 -684
rect 165 684 303 1116
rect 165 -1116 303 -684
rect 399 684 537 1116
rect 399 -1116 537 -684
rect 633 684 771 1116
rect 633 -1116 771 -684
rect 867 684 1005 1116
rect 867 -1116 1005 -684
rect 1101 684 1239 1116
rect 1101 -1116 1239 -684
rect 1335 684 1473 1116
rect 1335 -1116 1473 -684
rect 1569 684 1707 1116
rect 1569 -1116 1707 -684
rect 1803 684 1941 1116
rect 1803 -1116 1941 -684
rect 2037 684 2175 1116
rect 2037 -1116 2175 -684
rect 2271 684 2409 1116
rect 2271 -1116 2409 -684
rect 2505 684 2643 1116
rect 2505 -1116 2643 -684
rect 2739 684 2877 1116
rect 2739 -1116 2877 -684
rect 2973 684 3111 1116
rect 2973 -1116 3111 -684
<< xpolyres >>
rect -3111 -684 -2973 684
rect -2877 -684 -2739 684
rect -2643 -684 -2505 684
rect -2409 -684 -2271 684
rect -2175 -684 -2037 684
rect -1941 -684 -1803 684
rect -1707 -684 -1569 684
rect -1473 -684 -1335 684
rect -1239 -684 -1101 684
rect -1005 -684 -867 684
rect -771 -684 -633 684
rect -537 -684 -399 684
rect -303 -684 -165 684
rect -69 -684 69 684
rect 165 -684 303 684
rect 399 -684 537 684
rect 633 -684 771 684
rect 867 -684 1005 684
rect 1101 -684 1239 684
rect 1335 -684 1473 684
rect 1569 -684 1707 684
rect 1803 -684 1941 684
rect 2037 -684 2175 684
rect 2271 -684 2409 684
rect 2505 -684 2643 684
rect 2739 -684 2877 684
rect 2973 -684 3111 684
<< locali >>
rect -3241 1150 -3207 1166
rect 3207 1150 3241 1166
rect -3241 -1166 -3207 -1150
rect 3207 -1166 3241 -1150
rect -3161 -1246 -3145 -1212
rect 3145 -1246 3161 -1212
<< viali >>
rect -3095 701 -2989 1098
rect -2861 701 -2755 1098
rect -2627 701 -2521 1098
rect -2393 701 -2287 1098
rect -2159 701 -2053 1098
rect -1925 701 -1819 1098
rect -1691 701 -1585 1098
rect -1457 701 -1351 1098
rect -1223 701 -1117 1098
rect -989 701 -883 1098
rect -755 701 -649 1098
rect -521 701 -415 1098
rect -287 701 -181 1098
rect -53 701 53 1098
rect 181 701 287 1098
rect 415 701 521 1098
rect 649 701 755 1098
rect 883 701 989 1098
rect 1117 701 1223 1098
rect 1351 701 1457 1098
rect 1585 701 1691 1098
rect 1819 701 1925 1098
rect 2053 701 2159 1098
rect 2287 701 2393 1098
rect 2521 701 2627 1098
rect 2755 701 2861 1098
rect 2989 701 3095 1098
rect -3095 -1098 -2989 -701
rect -2861 -1098 -2755 -701
rect -2627 -1098 -2521 -701
rect -2393 -1098 -2287 -701
rect -2159 -1098 -2053 -701
rect -1925 -1098 -1819 -701
rect -1691 -1098 -1585 -701
rect -1457 -1098 -1351 -701
rect -1223 -1098 -1117 -701
rect -989 -1098 -883 -701
rect -755 -1098 -649 -701
rect -521 -1098 -415 -701
rect -287 -1098 -181 -701
rect -53 -1098 53 -701
rect 181 -1098 287 -701
rect 415 -1098 521 -701
rect 649 -1098 755 -701
rect 883 -1098 989 -701
rect 1117 -1098 1223 -701
rect 1351 -1098 1457 -701
rect 1585 -1098 1691 -701
rect 1819 -1098 1925 -701
rect 2053 -1098 2159 -701
rect 2287 -1098 2393 -701
rect 2521 -1098 2627 -701
rect 2755 -1098 2861 -701
rect 2989 -1098 3095 -701
<< metal1 >>
rect -3101 1098 -2983 1110
rect -3101 701 -3095 1098
rect -2989 701 -2983 1098
rect -3101 689 -2983 701
rect -2867 1098 -2749 1110
rect -2867 701 -2861 1098
rect -2755 701 -2749 1098
rect -2867 689 -2749 701
rect -2633 1098 -2515 1110
rect -2633 701 -2627 1098
rect -2521 701 -2515 1098
rect -2633 689 -2515 701
rect -2399 1098 -2281 1110
rect -2399 701 -2393 1098
rect -2287 701 -2281 1098
rect -2399 689 -2281 701
rect -2165 1098 -2047 1110
rect -2165 701 -2159 1098
rect -2053 701 -2047 1098
rect -2165 689 -2047 701
rect -1931 1098 -1813 1110
rect -1931 701 -1925 1098
rect -1819 701 -1813 1098
rect -1931 689 -1813 701
rect -1697 1098 -1579 1110
rect -1697 701 -1691 1098
rect -1585 701 -1579 1098
rect -1697 689 -1579 701
rect -1463 1098 -1345 1110
rect -1463 701 -1457 1098
rect -1351 701 -1345 1098
rect -1463 689 -1345 701
rect -1229 1098 -1111 1110
rect -1229 701 -1223 1098
rect -1117 701 -1111 1098
rect -1229 689 -1111 701
rect -995 1098 -877 1110
rect -995 701 -989 1098
rect -883 701 -877 1098
rect -995 689 -877 701
rect -761 1098 -643 1110
rect -761 701 -755 1098
rect -649 701 -643 1098
rect -761 689 -643 701
rect -527 1098 -409 1110
rect -527 701 -521 1098
rect -415 701 -409 1098
rect -527 689 -409 701
rect -293 1098 -175 1110
rect -293 701 -287 1098
rect -181 701 -175 1098
rect -293 689 -175 701
rect -59 1098 59 1110
rect -59 701 -53 1098
rect 53 701 59 1098
rect -59 689 59 701
rect 175 1098 293 1110
rect 175 701 181 1098
rect 287 701 293 1098
rect 175 689 293 701
rect 409 1098 527 1110
rect 409 701 415 1098
rect 521 701 527 1098
rect 409 689 527 701
rect 643 1098 761 1110
rect 643 701 649 1098
rect 755 701 761 1098
rect 643 689 761 701
rect 877 1098 995 1110
rect 877 701 883 1098
rect 989 701 995 1098
rect 877 689 995 701
rect 1111 1098 1229 1110
rect 1111 701 1117 1098
rect 1223 701 1229 1098
rect 1111 689 1229 701
rect 1345 1098 1463 1110
rect 1345 701 1351 1098
rect 1457 701 1463 1098
rect 1345 689 1463 701
rect 1579 1098 1697 1110
rect 1579 701 1585 1098
rect 1691 701 1697 1098
rect 1579 689 1697 701
rect 1813 1098 1931 1110
rect 1813 701 1819 1098
rect 1925 701 1931 1098
rect 1813 689 1931 701
rect 2047 1098 2165 1110
rect 2047 701 2053 1098
rect 2159 701 2165 1098
rect 2047 689 2165 701
rect 2281 1098 2399 1110
rect 2281 701 2287 1098
rect 2393 701 2399 1098
rect 2281 689 2399 701
rect 2515 1098 2633 1110
rect 2515 701 2521 1098
rect 2627 701 2633 1098
rect 2515 689 2633 701
rect 2749 1098 2867 1110
rect 2749 701 2755 1098
rect 2861 701 2867 1098
rect 2749 689 2867 701
rect 2983 1098 3101 1110
rect 2983 701 2989 1098
rect 3095 701 3101 1098
rect 2983 689 3101 701
rect -3101 -701 -2983 -689
rect -3101 -1098 -3095 -701
rect -2989 -1098 -2983 -701
rect -3101 -1110 -2983 -1098
rect -2867 -701 -2749 -689
rect -2867 -1098 -2861 -701
rect -2755 -1098 -2749 -701
rect -2867 -1110 -2749 -1098
rect -2633 -701 -2515 -689
rect -2633 -1098 -2627 -701
rect -2521 -1098 -2515 -701
rect -2633 -1110 -2515 -1098
rect -2399 -701 -2281 -689
rect -2399 -1098 -2393 -701
rect -2287 -1098 -2281 -701
rect -2399 -1110 -2281 -1098
rect -2165 -701 -2047 -689
rect -2165 -1098 -2159 -701
rect -2053 -1098 -2047 -701
rect -2165 -1110 -2047 -1098
rect -1931 -701 -1813 -689
rect -1931 -1098 -1925 -701
rect -1819 -1098 -1813 -701
rect -1931 -1110 -1813 -1098
rect -1697 -701 -1579 -689
rect -1697 -1098 -1691 -701
rect -1585 -1098 -1579 -701
rect -1697 -1110 -1579 -1098
rect -1463 -701 -1345 -689
rect -1463 -1098 -1457 -701
rect -1351 -1098 -1345 -701
rect -1463 -1110 -1345 -1098
rect -1229 -701 -1111 -689
rect -1229 -1098 -1223 -701
rect -1117 -1098 -1111 -701
rect -1229 -1110 -1111 -1098
rect -995 -701 -877 -689
rect -995 -1098 -989 -701
rect -883 -1098 -877 -701
rect -995 -1110 -877 -1098
rect -761 -701 -643 -689
rect -761 -1098 -755 -701
rect -649 -1098 -643 -701
rect -761 -1110 -643 -1098
rect -527 -701 -409 -689
rect -527 -1098 -521 -701
rect -415 -1098 -409 -701
rect -527 -1110 -409 -1098
rect -293 -701 -175 -689
rect -293 -1098 -287 -701
rect -181 -1098 -175 -701
rect -293 -1110 -175 -1098
rect -59 -701 59 -689
rect -59 -1098 -53 -701
rect 53 -1098 59 -701
rect -59 -1110 59 -1098
rect 175 -701 293 -689
rect 175 -1098 181 -701
rect 287 -1098 293 -701
rect 175 -1110 293 -1098
rect 409 -701 527 -689
rect 409 -1098 415 -701
rect 521 -1098 527 -701
rect 409 -1110 527 -1098
rect 643 -701 761 -689
rect 643 -1098 649 -701
rect 755 -1098 761 -701
rect 643 -1110 761 -1098
rect 877 -701 995 -689
rect 877 -1098 883 -701
rect 989 -1098 995 -701
rect 877 -1110 995 -1098
rect 1111 -701 1229 -689
rect 1111 -1098 1117 -701
rect 1223 -1098 1229 -701
rect 1111 -1110 1229 -1098
rect 1345 -701 1463 -689
rect 1345 -1098 1351 -701
rect 1457 -1098 1463 -701
rect 1345 -1110 1463 -1098
rect 1579 -701 1697 -689
rect 1579 -1098 1585 -701
rect 1691 -1098 1697 -701
rect 1579 -1110 1697 -1098
rect 1813 -701 1931 -689
rect 1813 -1098 1819 -701
rect 1925 -1098 1931 -701
rect 1813 -1110 1931 -1098
rect 2047 -701 2165 -689
rect 2047 -1098 2053 -701
rect 2159 -1098 2165 -701
rect 2047 -1110 2165 -1098
rect 2281 -701 2399 -689
rect 2281 -1098 2287 -701
rect 2393 -1098 2399 -701
rect 2281 -1110 2399 -1098
rect 2515 -701 2633 -689
rect 2515 -1098 2521 -701
rect 2627 -1098 2633 -701
rect 2515 -1110 2633 -1098
rect 2749 -701 2867 -689
rect 2749 -1098 2755 -701
rect 2861 -1098 2867 -701
rect 2749 -1110 2867 -1098
rect 2983 -701 3101 -689
rect 2983 -1098 2989 -701
rect 3095 -1098 3101 -701
rect 2983 -1110 3101 -1098
<< properties >>
string FIXED_BBOX -3224 -1229 3224 1229
string gencell sky130_fd_pr__res_xhigh_po_0p69
string library sky130
string parameters w 0.690 l 7.0 m 1 nx 27 wmin 0.690 lmin 0.50 rho 2000 val 20.835k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 0 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 0 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
