VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_cas_sensor_project
  CLASS BLOCK ;
  FOREIGN tt_um_cas_sensor_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 319.240 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    PORT
      LAYER met4 ;
        RECT 7.000 5.000 9.000 220.760 ;
    END
  END VAPWR
  OBS
      LAYER nwell ;
        RECT 35.000 154.745 109.440 156.350 ;
      LAYER pwell ;
        RECT 35.195 153.545 36.565 154.355 ;
        RECT 37.495 153.545 38.865 154.325 ;
        RECT 38.875 153.545 44.385 154.355 ;
        RECT 44.395 153.545 48.065 154.355 ;
        RECT 48.085 153.630 48.515 154.415 ;
        RECT 48.535 153.545 54.045 154.355 ;
        RECT 54.055 153.545 59.565 154.355 ;
        RECT 59.575 153.545 60.945 154.355 ;
        RECT 60.965 153.630 61.395 154.415 ;
        RECT 61.415 153.545 66.925 154.355 ;
        RECT 66.935 153.545 72.445 154.355 ;
        RECT 72.455 153.545 73.825 154.355 ;
        RECT 73.845 153.630 74.275 154.415 ;
        RECT 74.765 153.545 76.115 154.455 ;
        RECT 76.135 153.545 81.645 154.355 ;
        RECT 81.655 153.545 85.325 154.355 ;
        RECT 85.335 153.545 86.705 154.355 ;
        RECT 86.725 153.630 87.155 154.415 ;
        RECT 87.175 153.545 92.685 154.355 ;
        RECT 92.695 153.545 98.205 154.355 ;
        RECT 98.215 153.545 99.585 154.355 ;
        RECT 99.605 153.630 100.035 154.415 ;
        RECT 100.055 153.545 105.565 154.355 ;
        RECT 105.575 153.545 107.405 154.355 ;
        RECT 107.875 153.545 109.245 154.355 ;
        RECT 35.335 153.335 35.505 153.545 ;
        RECT 36.715 153.335 36.885 153.525 ;
        RECT 37.645 153.355 37.815 153.545 ;
        RECT 39.015 153.355 39.185 153.545 ;
        RECT 42.235 153.335 42.405 153.525 ;
        RECT 44.535 153.355 44.705 153.545 ;
        RECT 47.755 153.335 47.925 153.525 ;
        RECT 48.675 153.355 48.845 153.545 ;
        RECT 53.275 153.335 53.445 153.525 ;
        RECT 54.195 153.355 54.365 153.545 ;
        RECT 55.110 153.385 55.230 153.495 ;
        RECT 55.580 153.335 55.750 153.525 ;
        RECT 59.255 153.335 59.425 153.525 ;
        RECT 59.715 153.335 59.885 153.545 ;
        RECT 61.555 153.355 61.725 153.545 ;
        RECT 62.475 153.335 62.645 153.525 ;
        RECT 63.855 153.335 64.025 153.525 ;
        RECT 64.310 153.385 64.430 153.495 ;
        RECT 64.775 153.335 64.945 153.525 ;
        RECT 66.155 153.335 66.325 153.525 ;
        RECT 67.075 153.355 67.245 153.545 ;
        RECT 72.595 153.355 72.765 153.545 ;
        RECT 74.430 153.385 74.550 153.495 ;
        RECT 74.895 153.355 75.065 153.545 ;
        RECT 75.365 153.380 75.525 153.490 ;
        RECT 76.275 153.335 76.445 153.545 ;
        RECT 81.795 153.355 81.965 153.545 ;
        RECT 85.475 153.355 85.645 153.545 ;
        RECT 86.395 153.335 86.565 153.525 ;
        RECT 87.315 153.335 87.485 153.545 ;
        RECT 92.835 153.355 93.005 153.545 ;
        RECT 96.515 153.335 96.685 153.525 ;
        RECT 97.895 153.335 98.065 153.525 ;
        RECT 98.355 153.355 98.525 153.545 ;
        RECT 100.195 153.355 100.365 153.545 ;
        RECT 103.415 153.335 103.585 153.525 ;
        RECT 105.715 153.355 105.885 153.545 ;
        RECT 107.105 153.380 107.265 153.490 ;
        RECT 107.550 153.385 107.670 153.495 ;
        RECT 108.935 153.335 109.105 153.545 ;
        RECT 35.195 152.525 36.565 153.335 ;
        RECT 36.575 152.525 42.085 153.335 ;
        RECT 42.095 152.525 47.605 153.335 ;
        RECT 47.615 152.525 53.125 153.335 ;
        RECT 53.135 152.525 54.965 153.335 ;
        RECT 55.435 152.425 58.045 153.335 ;
        RECT 58.205 152.425 59.555 153.335 ;
        RECT 59.575 152.525 60.945 153.335 ;
        RECT 60.965 152.465 61.395 153.250 ;
        RECT 61.425 152.425 62.775 153.335 ;
        RECT 62.805 152.425 64.155 153.335 ;
        RECT 64.645 152.425 65.995 153.335 ;
        RECT 66.015 152.655 75.205 153.335 ;
        RECT 76.135 152.655 85.325 153.335 ;
        RECT 70.525 152.435 71.455 152.655 ;
        RECT 74.285 152.425 75.205 152.655 ;
        RECT 80.645 152.435 81.575 152.655 ;
        RECT 84.405 152.425 85.325 152.655 ;
        RECT 85.345 152.425 86.695 153.335 ;
        RECT 86.725 152.465 87.155 153.250 ;
        RECT 87.175 152.655 96.365 153.335 ;
        RECT 91.685 152.435 92.615 152.655 ;
        RECT 95.445 152.425 96.365 152.655 ;
        RECT 96.385 152.425 97.735 153.335 ;
        RECT 97.755 152.525 103.265 153.335 ;
        RECT 103.275 152.525 106.945 153.335 ;
        RECT 107.875 152.525 109.245 153.335 ;
      LAYER nwell ;
        RECT 35.000 149.305 109.440 152.135 ;
      LAYER pwell ;
        RECT 35.195 148.105 36.565 148.915 ;
        RECT 36.575 148.105 42.085 148.915 ;
        RECT 42.095 148.105 47.605 148.915 ;
        RECT 48.085 148.190 48.515 148.975 ;
        RECT 48.535 148.105 54.045 148.915 ;
        RECT 54.055 148.105 55.425 148.915 ;
        RECT 59.945 148.785 60.875 149.005 ;
        RECT 63.705 148.785 64.625 149.015 ;
        RECT 67.290 148.785 68.210 149.015 ;
        RECT 55.435 148.105 64.625 148.785 ;
        RECT 64.745 148.105 68.210 148.785 ;
        RECT 68.315 148.105 71.065 149.015 ;
        RECT 71.085 148.105 72.435 149.015 ;
        RECT 72.455 148.105 73.825 148.915 ;
        RECT 73.845 148.190 74.275 148.975 ;
        RECT 74.390 148.785 75.310 149.015 ;
        RECT 78.460 148.785 79.805 149.015 ;
        RECT 74.390 148.105 77.855 148.785 ;
        RECT 77.975 148.105 79.805 148.785 ;
        RECT 79.815 148.105 83.485 148.915 ;
        RECT 83.965 148.105 85.315 149.015 ;
        RECT 85.795 148.105 87.625 149.015 ;
        RECT 87.635 148.105 90.385 148.915 ;
        RECT 90.865 148.105 92.215 149.015 ;
        RECT 92.235 148.105 97.745 148.915 ;
        RECT 97.755 148.105 99.585 148.915 ;
        RECT 99.605 148.190 100.035 148.975 ;
        RECT 100.055 148.105 105.565 148.915 ;
        RECT 105.575 148.105 107.405 148.915 ;
        RECT 107.875 148.105 109.245 148.915 ;
        RECT 35.335 147.895 35.505 148.105 ;
        RECT 36.715 147.895 36.885 148.105 ;
        RECT 42.235 147.895 42.405 148.105 ;
        RECT 47.755 148.055 47.925 148.085 ;
        RECT 47.750 147.945 47.925 148.055 ;
        RECT 47.755 147.915 47.925 147.945 ;
        RECT 48.675 147.915 48.845 148.105 ;
        RECT 49.135 147.895 49.305 148.085 ;
        RECT 51.895 147.895 52.065 148.085 ;
        RECT 52.355 147.895 52.525 148.085 ;
        RECT 54.195 147.915 54.365 148.105 ;
        RECT 55.575 147.915 55.745 148.105 ;
        RECT 56.030 147.945 56.150 148.055 ;
        RECT 58.335 147.895 58.505 148.085 ;
        RECT 35.195 147.085 36.565 147.895 ;
        RECT 36.575 147.085 42.085 147.895 ;
        RECT 42.095 147.085 47.605 147.895 ;
        RECT 48.995 147.085 50.825 147.895 ;
        RECT 50.845 146.985 52.195 147.895 ;
        RECT 52.215 147.085 55.885 147.895 ;
        RECT 56.355 146.985 58.645 147.895 ;
        RECT 58.655 147.865 59.610 147.895 ;
        RECT 60.640 147.865 60.810 148.085 ;
        RECT 61.565 147.940 61.725 148.050 ;
        RECT 62.475 147.895 62.645 148.085 ;
        RECT 64.775 147.915 64.945 148.105 ;
        RECT 58.655 147.185 60.935 147.865 ;
        RECT 58.655 146.985 59.610 147.185 ;
        RECT 60.965 147.025 61.395 147.810 ;
        RECT 62.445 147.215 65.910 147.895 ;
        RECT 64.990 146.985 65.910 147.215 ;
        RECT 66.015 147.865 66.970 147.895 ;
        RECT 68.000 147.865 68.170 148.085 ;
        RECT 68.450 147.915 68.620 148.085 ;
        RECT 70.755 147.915 70.925 148.105 ;
        RECT 71.215 147.915 71.385 148.105 ;
        RECT 72.595 147.915 72.765 148.105 ;
        RECT 68.485 147.895 68.620 147.915 ;
        RECT 66.015 147.185 68.295 147.865 ;
        RECT 66.015 146.985 66.970 147.185 ;
        RECT 68.485 146.985 71.985 147.895 ;
        RECT 71.995 147.865 72.930 147.895 ;
        RECT 74.890 147.865 75.060 148.085 ;
        RECT 76.280 147.895 76.450 148.085 ;
        RECT 76.730 147.915 76.900 148.085 ;
        RECT 77.655 147.915 77.825 148.105 ;
        RECT 78.115 147.915 78.285 148.105 ;
        RECT 79.955 147.915 80.125 148.105 ;
        RECT 80.410 147.945 80.530 148.055 ;
        RECT 76.765 147.895 76.900 147.915 ;
        RECT 71.995 147.665 75.060 147.865 ;
        RECT 71.995 147.185 75.205 147.665 ;
        RECT 71.995 146.985 72.945 147.185 ;
        RECT 74.275 146.985 75.205 147.185 ;
        RECT 75.215 146.985 76.565 147.895 ;
        RECT 76.765 146.985 80.265 147.895 ;
        RECT 80.870 147.865 81.040 148.085 ;
        RECT 83.180 147.895 83.350 148.085 ;
        RECT 83.630 147.945 83.750 148.055 ;
        RECT 85.015 147.915 85.185 148.105 ;
        RECT 85.940 148.085 86.110 148.105 ;
        RECT 85.470 147.945 85.590 148.055 ;
        RECT 85.930 147.915 86.110 148.085 ;
        RECT 86.390 147.945 86.510 148.055 ;
        RECT 85.930 147.895 86.100 147.915 ;
        RECT 87.315 147.895 87.485 148.085 ;
        RECT 87.775 147.915 87.945 148.105 ;
        RECT 90.535 148.055 90.705 148.085 ;
        RECT 90.530 147.945 90.705 148.055 ;
        RECT 90.535 147.895 90.705 147.945 ;
        RECT 90.995 147.915 91.165 148.105 ;
        RECT 92.375 147.915 92.545 148.105 ;
        RECT 96.055 147.895 96.225 148.085 ;
        RECT 97.895 147.915 98.065 148.105 ;
        RECT 100.195 147.915 100.365 148.105 ;
        RECT 101.575 147.895 101.745 148.085 ;
        RECT 105.715 147.915 105.885 148.105 ;
        RECT 107.105 147.940 107.265 148.050 ;
        RECT 107.550 147.945 107.670 148.055 ;
        RECT 108.935 147.895 109.105 148.105 ;
        RECT 82.070 147.865 83.025 147.895 ;
        RECT 80.745 147.185 83.025 147.865 ;
        RECT 82.070 146.985 83.025 147.185 ;
        RECT 83.035 146.985 84.865 147.895 ;
        RECT 84.895 146.985 86.245 147.895 ;
        RECT 86.725 147.025 87.155 147.810 ;
        RECT 87.175 146.985 90.385 147.895 ;
        RECT 90.395 147.085 95.905 147.895 ;
        RECT 95.915 147.085 101.425 147.895 ;
        RECT 101.435 147.085 106.945 147.895 ;
        RECT 107.875 147.085 109.245 147.895 ;
      LAYER nwell ;
        RECT 35.000 143.865 109.440 146.695 ;
      LAYER pwell ;
        RECT 35.195 142.665 36.565 143.475 ;
        RECT 36.575 142.665 42.085 143.475 ;
        RECT 42.095 142.665 47.605 143.475 ;
        RECT 48.085 142.750 48.515 143.535 ;
        RECT 48.535 142.665 54.045 143.475 ;
        RECT 55.060 142.665 64.165 143.345 ;
        RECT 64.635 142.665 73.740 143.345 ;
        RECT 73.845 142.750 74.275 143.535 ;
        RECT 74.295 142.895 77.495 143.575 ;
        RECT 74.440 142.665 77.495 142.895 ;
        RECT 77.515 142.665 81.185 143.475 ;
        RECT 82.125 142.665 83.475 143.575 ;
        RECT 83.495 142.665 89.005 143.475 ;
        RECT 89.015 142.665 94.525 143.475 ;
        RECT 94.535 142.665 95.905 143.475 ;
        RECT 95.925 142.665 97.275 143.575 ;
        RECT 97.295 142.665 99.125 143.475 ;
        RECT 99.605 142.750 100.035 143.535 ;
        RECT 100.055 142.665 105.565 143.475 ;
        RECT 105.575 142.665 107.405 143.475 ;
        RECT 107.875 142.665 109.245 143.475 ;
        RECT 35.335 142.455 35.505 142.665 ;
        RECT 36.715 142.455 36.885 142.665 ;
        RECT 42.235 142.615 42.405 142.665 ;
        RECT 42.230 142.505 42.405 142.615 ;
        RECT 42.235 142.475 42.405 142.505 ;
        RECT 42.695 142.455 42.865 142.645 ;
        RECT 47.750 142.505 47.870 142.615 ;
        RECT 48.675 142.475 48.845 142.665 ;
        RECT 51.895 142.455 52.065 142.645 ;
        RECT 54.205 142.510 54.365 142.620 ;
        RECT 61.560 142.455 61.730 142.645 ;
        RECT 63.855 142.475 64.025 142.665 ;
        RECT 64.310 142.505 64.430 142.615 ;
        RECT 64.775 142.475 64.945 142.665 ;
        RECT 65.245 142.500 65.405 142.610 ;
        RECT 67.080 142.455 67.250 142.645 ;
        RECT 67.535 142.455 67.705 142.645 ;
        RECT 35.195 141.645 36.565 142.455 ;
        RECT 36.575 141.645 42.085 142.455 ;
        RECT 42.555 141.775 51.745 142.455 ;
        RECT 51.755 141.775 60.945 142.455 ;
        RECT 47.065 141.555 47.995 141.775 ;
        RECT 50.825 141.545 51.745 141.775 ;
        RECT 56.265 141.555 57.195 141.775 ;
        RECT 60.025 141.545 60.945 141.775 ;
        RECT 60.965 141.585 61.395 142.370 ;
        RECT 61.415 141.775 65.000 142.455 ;
        RECT 61.415 141.545 62.335 141.775 ;
        RECT 66.015 141.545 67.365 142.455 ;
        RECT 67.395 141.645 71.065 142.455 ;
        RECT 71.220 142.425 71.390 142.645 ;
        RECT 74.440 142.475 74.610 142.665 ;
        RECT 74.890 142.455 75.060 142.645 ;
        RECT 75.350 142.505 75.470 142.615 ;
        RECT 75.815 142.455 75.985 142.645 ;
        RECT 77.195 142.455 77.365 142.645 ;
        RECT 77.655 142.475 77.825 142.665 ;
        RECT 72.880 142.425 73.825 142.455 ;
        RECT 71.075 141.745 73.825 142.425 ;
        RECT 72.880 141.545 73.825 141.745 ;
        RECT 73.855 141.545 75.205 142.455 ;
        RECT 75.685 141.545 77.035 142.455 ;
        RECT 77.055 141.645 78.425 142.455 ;
        RECT 78.575 142.425 78.745 142.645 ;
        RECT 81.345 142.510 81.505 142.620 ;
        RECT 81.805 142.500 81.965 142.610 ;
        RECT 82.255 142.475 82.425 142.665 ;
        RECT 83.635 142.475 83.805 142.665 ;
        RECT 85.930 142.455 86.100 142.645 ;
        RECT 86.390 142.505 86.510 142.615 ;
        RECT 87.315 142.455 87.485 142.645 ;
        RECT 89.155 142.475 89.325 142.665 ;
        RECT 94.675 142.475 94.845 142.665 ;
        RECT 96.055 142.475 96.225 142.665 ;
        RECT 96.515 142.455 96.685 142.645 ;
        RECT 97.435 142.475 97.605 142.665 ;
        RECT 99.270 142.505 99.390 142.615 ;
        RECT 100.195 142.475 100.365 142.665 ;
        RECT 102.035 142.455 102.205 142.645 ;
        RECT 105.715 142.475 105.885 142.665 ;
        RECT 107.550 142.505 107.670 142.615 ;
        RECT 108.935 142.455 109.105 142.665 ;
        RECT 80.700 142.425 81.645 142.455 ;
        RECT 78.575 142.225 81.645 142.425 ;
        RECT 78.435 141.745 81.645 142.225 ;
        RECT 78.435 141.545 79.365 141.745 ;
        RECT 80.700 141.545 81.645 141.745 ;
        RECT 82.575 141.545 86.245 142.455 ;
        RECT 86.725 141.585 87.155 142.370 ;
        RECT 87.175 141.775 96.365 142.455 ;
        RECT 91.685 141.555 92.615 141.775 ;
        RECT 95.445 141.545 96.365 141.775 ;
        RECT 96.375 141.645 101.885 142.455 ;
        RECT 101.895 141.645 107.405 142.455 ;
        RECT 107.875 141.645 109.245 142.455 ;
      LAYER nwell ;
        RECT 35.000 138.425 109.440 141.255 ;
      LAYER pwell ;
        RECT 35.195 137.225 36.565 138.035 ;
        RECT 36.575 137.225 42.085 138.035 ;
        RECT 42.095 137.225 47.605 138.035 ;
        RECT 48.085 137.310 48.515 138.095 ;
        RECT 48.535 137.225 54.045 138.035 ;
        RECT 54.055 137.225 55.425 138.035 ;
        RECT 55.445 137.225 56.795 138.135 ;
        RECT 56.815 137.225 58.645 138.035 ;
        RECT 59.195 137.225 62.195 138.135 ;
        RECT 62.335 137.225 66.005 138.135 ;
        RECT 66.110 137.905 67.030 138.135 ;
        RECT 66.110 137.225 69.575 137.905 ;
        RECT 70.150 137.455 71.985 138.135 ;
        RECT 70.150 137.225 71.840 137.455 ;
        RECT 71.995 137.225 73.825 138.035 ;
        RECT 73.845 137.310 74.275 138.095 ;
        RECT 74.295 137.225 75.665 138.035 ;
        RECT 75.695 137.225 77.045 138.135 ;
        RECT 77.055 137.455 80.255 138.135 ;
        RECT 89.570 137.905 90.490 138.135 ;
        RECT 77.200 137.225 80.255 137.455 ;
        RECT 80.275 137.225 89.380 137.905 ;
        RECT 89.570 137.225 93.035 137.905 ;
        RECT 93.155 137.225 94.985 138.135 ;
        RECT 95.005 137.225 96.355 138.135 ;
        RECT 96.375 137.225 99.125 138.035 ;
        RECT 99.605 137.310 100.035 138.095 ;
        RECT 100.055 137.225 103.725 138.035 ;
        RECT 104.665 137.225 106.015 138.135 ;
        RECT 106.035 137.225 107.865 138.035 ;
        RECT 107.875 137.225 109.245 138.035 ;
        RECT 35.335 137.015 35.505 137.225 ;
        RECT 36.715 137.015 36.885 137.225 ;
        RECT 42.235 137.015 42.405 137.225 ;
        RECT 47.755 137.175 47.925 137.205 ;
        RECT 47.750 137.065 47.925 137.175 ;
        RECT 47.755 137.015 47.925 137.065 ;
        RECT 48.675 137.035 48.845 137.225 ;
        RECT 51.430 137.065 51.550 137.175 ;
        RECT 51.895 137.015 52.065 137.205 ;
        RECT 54.195 137.035 54.365 137.225 ;
        RECT 55.575 137.035 55.745 137.225 ;
        RECT 56.955 137.035 57.125 137.225 ;
        RECT 58.790 137.065 58.910 137.175 ;
        RECT 59.255 137.035 59.425 137.225 ;
        RECT 62.480 137.205 62.650 137.225 ;
        RECT 62.475 137.035 62.650 137.205 ;
        RECT 62.475 137.015 62.645 137.035 ;
        RECT 62.935 137.015 63.105 137.205 ;
        RECT 65.690 137.065 65.810 137.175 ;
        RECT 66.155 137.015 66.325 137.205 ;
        RECT 67.535 137.015 67.705 137.205 ;
        RECT 69.375 137.035 69.545 137.225 ;
        RECT 70.295 137.015 70.465 137.205 ;
        RECT 71.670 137.035 71.840 137.225 ;
        RECT 72.135 137.035 72.305 137.225 ;
        RECT 74.435 137.035 74.605 137.225 ;
        RECT 76.275 137.015 76.445 137.205 ;
        RECT 76.730 137.170 76.900 137.225 ;
        RECT 76.730 137.060 76.905 137.170 ;
        RECT 76.730 137.035 76.900 137.060 ;
        RECT 77.200 137.035 77.370 137.225 ;
        RECT 77.660 137.015 77.830 137.205 ;
        RECT 35.195 136.205 36.565 137.015 ;
        RECT 36.575 136.205 42.085 137.015 ;
        RECT 42.095 136.205 47.605 137.015 ;
        RECT 47.615 136.205 51.285 137.015 ;
        RECT 51.755 136.335 60.945 137.015 ;
        RECT 56.265 136.115 57.195 136.335 ;
        RECT 60.025 136.105 60.945 136.335 ;
        RECT 60.965 136.145 61.395 136.930 ;
        RECT 61.425 136.105 62.775 137.015 ;
        RECT 62.795 136.205 65.545 137.015 ;
        RECT 66.025 136.105 67.375 137.015 ;
        RECT 67.395 136.205 70.145 137.015 ;
        RECT 70.265 136.335 73.730 137.015 ;
        RECT 72.810 136.105 73.730 136.335 ;
        RECT 73.845 136.105 76.575 137.015 ;
        RECT 77.515 136.105 79.345 137.015 ;
        RECT 79.500 136.985 79.670 137.205 ;
        RECT 80.415 137.035 80.585 137.225 ;
        RECT 85.470 137.015 85.640 137.205 ;
        RECT 85.945 137.060 86.105 137.170 ;
        RECT 87.315 137.015 87.485 137.205 ;
        RECT 92.835 137.035 93.005 137.225 ;
        RECT 93.300 137.035 93.470 137.225 ;
        RECT 95.135 137.035 95.305 137.225 ;
        RECT 96.515 137.015 96.685 137.225 ;
        RECT 99.270 137.065 99.390 137.175 ;
        RECT 100.195 137.035 100.365 137.225 ;
        RECT 102.035 137.015 102.205 137.205 ;
        RECT 103.885 137.070 104.045 137.180 ;
        RECT 104.795 137.035 104.965 137.225 ;
        RECT 106.175 137.035 106.345 137.225 ;
        RECT 107.550 137.065 107.670 137.175 ;
        RECT 108.935 137.015 109.105 137.225 ;
        RECT 81.160 136.985 82.105 137.015 ;
        RECT 79.355 136.305 82.105 136.985 ;
        RECT 81.160 136.105 82.105 136.305 ;
        RECT 82.115 136.105 85.785 137.015 ;
        RECT 86.725 136.145 87.155 136.930 ;
        RECT 87.175 136.335 96.365 137.015 ;
        RECT 91.685 136.115 92.615 136.335 ;
        RECT 95.445 136.105 96.365 136.335 ;
        RECT 96.375 136.205 101.885 137.015 ;
        RECT 101.895 136.205 107.405 137.015 ;
        RECT 107.875 136.205 109.245 137.015 ;
      LAYER nwell ;
        RECT 35.000 132.985 109.440 135.815 ;
      LAYER pwell ;
        RECT 35.195 131.785 36.565 132.595 ;
        RECT 36.575 131.785 42.085 132.595 ;
        RECT 42.095 131.785 47.605 132.595 ;
        RECT 48.085 131.870 48.515 132.655 ;
        RECT 48.535 131.785 54.045 132.595 ;
        RECT 54.055 131.785 59.565 132.595 ;
        RECT 59.575 131.785 61.405 132.595 ;
        RECT 62.775 132.465 63.695 132.685 ;
        RECT 69.775 132.585 70.695 132.695 ;
        RECT 68.360 132.465 70.695 132.585 ;
        RECT 61.415 131.785 70.695 132.465 ;
        RECT 71.075 131.785 72.445 132.595 ;
        RECT 72.465 131.785 73.815 132.695 ;
        RECT 73.845 131.870 74.275 132.655 ;
        RECT 74.390 132.465 75.310 132.695 ;
        RECT 79.335 132.465 80.255 132.685 ;
        RECT 85.850 132.585 87.620 132.695 ;
        RECT 84.920 132.465 87.620 132.585 ;
        RECT 74.390 131.785 77.855 132.465 ;
        RECT 77.975 131.785 87.620 132.465 ;
        RECT 87.635 131.785 89.465 132.595 ;
        RECT 89.485 131.785 90.835 132.695 ;
        RECT 90.855 131.785 96.365 132.595 ;
        RECT 96.375 131.785 99.125 132.595 ;
        RECT 99.605 131.870 100.035 132.655 ;
        RECT 100.055 131.785 105.565 132.595 ;
        RECT 105.575 131.785 107.405 132.595 ;
        RECT 107.875 131.785 109.245 132.595 ;
        RECT 35.335 131.575 35.505 131.785 ;
        RECT 36.715 131.575 36.885 131.785 ;
        RECT 42.235 131.575 42.405 131.785 ;
        RECT 47.755 131.735 47.925 131.765 ;
        RECT 47.750 131.625 47.925 131.735 ;
        RECT 47.755 131.575 47.925 131.625 ;
        RECT 48.675 131.595 48.845 131.785 ;
        RECT 53.275 131.575 53.445 131.765 ;
        RECT 54.195 131.595 54.365 131.785 ;
        RECT 58.795 131.575 58.965 131.765 ;
        RECT 59.715 131.595 59.885 131.785 ;
        RECT 60.630 131.625 60.750 131.735 ;
        RECT 61.555 131.575 61.725 131.785 ;
        RECT 63.390 131.625 63.510 131.735 ;
        RECT 67.075 131.575 67.245 131.765 ;
        RECT 67.535 131.575 67.705 131.765 ;
        RECT 71.215 131.595 71.385 131.785 ;
        RECT 73.515 131.595 73.685 131.785 ;
        RECT 77.655 131.595 77.825 131.785 ;
        RECT 78.115 131.575 78.285 131.785 ;
        RECT 78.575 131.575 78.745 131.765 ;
        RECT 82.265 131.620 82.425 131.730 ;
        RECT 84.095 131.575 84.265 131.765 ;
        RECT 84.555 131.575 84.725 131.765 ;
        RECT 86.390 131.625 86.510 131.735 ;
        RECT 87.315 131.575 87.485 131.765 ;
        RECT 87.775 131.595 87.945 131.785 ;
        RECT 89.615 131.595 89.785 131.785 ;
        RECT 90.995 131.595 91.165 131.785 ;
        RECT 92.835 131.575 93.005 131.765 ;
        RECT 96.515 131.595 96.685 131.785 ;
        RECT 98.355 131.575 98.525 131.765 ;
        RECT 99.270 131.625 99.390 131.735 ;
        RECT 100.195 131.595 100.365 131.785 ;
        RECT 103.875 131.575 104.045 131.765 ;
        RECT 105.715 131.595 105.885 131.785 ;
        RECT 107.550 131.625 107.670 131.735 ;
        RECT 108.935 131.575 109.105 131.785 ;
        RECT 35.195 130.765 36.565 131.575 ;
        RECT 36.575 130.765 42.085 131.575 ;
        RECT 42.095 130.765 47.605 131.575 ;
        RECT 47.615 130.765 53.125 131.575 ;
        RECT 53.135 130.765 58.645 131.575 ;
        RECT 58.655 130.765 60.485 131.575 ;
        RECT 60.965 130.705 61.395 131.490 ;
        RECT 61.415 130.765 63.245 131.575 ;
        RECT 63.810 130.895 67.275 131.575 ;
        RECT 63.810 130.665 64.730 130.895 ;
        RECT 67.395 130.765 68.765 131.575 ;
        RECT 68.780 130.895 78.425 131.575 ;
        RECT 68.780 130.775 71.480 130.895 ;
        RECT 68.780 130.665 70.550 130.775 ;
        RECT 76.145 130.675 77.065 130.895 ;
        RECT 78.435 130.765 82.105 131.575 ;
        RECT 83.045 130.665 84.395 131.575 ;
        RECT 84.415 130.765 86.245 131.575 ;
        RECT 86.725 130.705 87.155 131.490 ;
        RECT 87.175 130.765 92.685 131.575 ;
        RECT 92.695 130.765 98.205 131.575 ;
        RECT 98.215 130.765 103.725 131.575 ;
        RECT 103.735 130.765 107.405 131.575 ;
        RECT 107.875 130.765 109.245 131.575 ;
      LAYER nwell ;
        RECT 35.000 127.545 109.440 130.375 ;
      LAYER pwell ;
        RECT 35.195 126.345 36.565 127.155 ;
        RECT 36.575 126.345 42.085 127.155 ;
        RECT 42.095 126.345 47.605 127.155 ;
        RECT 48.085 126.430 48.515 127.215 ;
        RECT 48.535 126.345 54.045 127.155 ;
        RECT 54.055 126.345 59.565 127.155 ;
        RECT 59.575 126.345 63.245 127.155 ;
        RECT 63.715 126.345 66.465 127.255 ;
        RECT 66.475 126.345 71.985 127.155 ;
        RECT 71.995 126.345 73.825 127.155 ;
        RECT 73.845 126.430 74.275 127.215 ;
        RECT 74.295 126.345 79.805 127.155 ;
        RECT 79.815 126.345 85.325 127.155 ;
        RECT 85.335 126.345 90.845 127.155 ;
        RECT 90.855 126.345 96.365 127.155 ;
        RECT 96.375 126.345 99.125 127.155 ;
        RECT 99.605 126.430 100.035 127.215 ;
        RECT 100.055 126.345 105.565 127.155 ;
        RECT 105.575 126.345 107.405 127.155 ;
        RECT 107.875 126.345 109.245 127.155 ;
        RECT 35.335 126.135 35.505 126.345 ;
        RECT 36.715 126.135 36.885 126.345 ;
        RECT 42.235 126.135 42.405 126.345 ;
        RECT 47.755 126.295 47.925 126.325 ;
        RECT 47.750 126.185 47.925 126.295 ;
        RECT 47.755 126.135 47.925 126.185 ;
        RECT 48.675 126.155 48.845 126.345 ;
        RECT 53.275 126.135 53.445 126.325 ;
        RECT 54.195 126.155 54.365 126.345 ;
        RECT 58.795 126.135 58.965 126.325 ;
        RECT 59.715 126.155 59.885 126.345 ;
        RECT 60.630 126.185 60.750 126.295 ;
        RECT 61.555 126.135 61.725 126.325 ;
        RECT 63.390 126.185 63.510 126.295 ;
        RECT 63.855 126.155 64.025 126.345 ;
        RECT 66.615 126.155 66.785 126.345 ;
        RECT 67.075 126.135 67.245 126.325 ;
        RECT 72.135 126.155 72.305 126.345 ;
        RECT 72.595 126.135 72.765 126.325 ;
        RECT 74.435 126.155 74.605 126.345 ;
        RECT 78.115 126.135 78.285 126.325 ;
        RECT 79.955 126.155 80.125 126.345 ;
        RECT 83.635 126.135 83.805 126.325 ;
        RECT 85.475 126.155 85.645 126.345 ;
        RECT 86.390 126.185 86.510 126.295 ;
        RECT 87.315 126.135 87.485 126.325 ;
        RECT 90.995 126.155 91.165 126.345 ;
        RECT 92.835 126.135 93.005 126.325 ;
        RECT 96.515 126.155 96.685 126.345 ;
        RECT 98.355 126.135 98.525 126.325 ;
        RECT 99.270 126.185 99.390 126.295 ;
        RECT 100.195 126.155 100.365 126.345 ;
        RECT 103.875 126.135 104.045 126.325 ;
        RECT 105.715 126.155 105.885 126.345 ;
        RECT 107.550 126.185 107.670 126.295 ;
        RECT 108.935 126.135 109.105 126.345 ;
        RECT 35.195 125.325 36.565 126.135 ;
        RECT 36.575 125.325 42.085 126.135 ;
        RECT 42.095 125.325 47.605 126.135 ;
        RECT 47.615 125.325 53.125 126.135 ;
        RECT 53.135 125.325 58.645 126.135 ;
        RECT 58.655 125.325 60.485 126.135 ;
        RECT 60.965 125.265 61.395 126.050 ;
        RECT 61.415 125.325 66.925 126.135 ;
        RECT 66.935 125.325 72.445 126.135 ;
        RECT 72.455 125.325 77.965 126.135 ;
        RECT 77.975 125.325 83.485 126.135 ;
        RECT 83.495 125.325 86.245 126.135 ;
        RECT 86.725 125.265 87.155 126.050 ;
        RECT 87.175 125.325 92.685 126.135 ;
        RECT 92.695 125.325 98.205 126.135 ;
        RECT 98.215 125.325 103.725 126.135 ;
        RECT 103.735 125.325 107.405 126.135 ;
        RECT 107.875 125.325 109.245 126.135 ;
      LAYER nwell ;
        RECT 35.000 122.105 109.440 124.935 ;
      LAYER pwell ;
        RECT 35.195 120.905 36.565 121.715 ;
        RECT 36.575 120.905 42.085 121.715 ;
        RECT 42.095 120.905 47.605 121.715 ;
        RECT 48.085 120.990 48.515 121.775 ;
        RECT 48.535 120.905 54.045 121.715 ;
        RECT 54.055 120.905 59.565 121.715 ;
        RECT 59.575 120.905 65.085 121.715 ;
        RECT 65.095 120.905 70.605 121.715 ;
        RECT 70.615 120.905 73.365 121.715 ;
        RECT 73.845 120.990 74.275 121.775 ;
        RECT 74.295 120.905 79.805 121.715 ;
        RECT 79.815 120.905 85.325 121.715 ;
        RECT 85.335 120.905 90.845 121.715 ;
        RECT 90.855 120.905 96.365 121.715 ;
        RECT 96.375 120.905 99.125 121.715 ;
        RECT 99.605 120.990 100.035 121.775 ;
        RECT 100.055 120.905 105.565 121.715 ;
        RECT 105.575 120.905 107.405 121.715 ;
        RECT 107.875 120.905 109.245 121.715 ;
        RECT 35.335 120.695 35.505 120.905 ;
        RECT 36.715 120.695 36.885 120.905 ;
        RECT 42.235 120.695 42.405 120.905 ;
        RECT 47.755 120.855 47.925 120.885 ;
        RECT 47.750 120.745 47.925 120.855 ;
        RECT 47.755 120.695 47.925 120.745 ;
        RECT 48.675 120.715 48.845 120.905 ;
        RECT 53.275 120.695 53.445 120.885 ;
        RECT 54.195 120.715 54.365 120.905 ;
        RECT 58.795 120.695 58.965 120.885 ;
        RECT 59.715 120.715 59.885 120.905 ;
        RECT 60.630 120.745 60.750 120.855 ;
        RECT 61.555 120.695 61.725 120.885 ;
        RECT 65.235 120.715 65.405 120.905 ;
        RECT 67.075 120.695 67.245 120.885 ;
        RECT 70.755 120.715 70.925 120.905 ;
        RECT 72.595 120.695 72.765 120.885 ;
        RECT 73.510 120.745 73.630 120.855 ;
        RECT 74.435 120.715 74.605 120.905 ;
        RECT 78.115 120.695 78.285 120.885 ;
        RECT 79.955 120.715 80.125 120.905 ;
        RECT 83.635 120.695 83.805 120.885 ;
        RECT 85.475 120.715 85.645 120.905 ;
        RECT 86.390 120.745 86.510 120.855 ;
        RECT 87.315 120.695 87.485 120.885 ;
        RECT 90.995 120.715 91.165 120.905 ;
        RECT 92.835 120.695 93.005 120.885 ;
        RECT 96.515 120.715 96.685 120.905 ;
        RECT 98.355 120.695 98.525 120.885 ;
        RECT 99.270 120.745 99.390 120.855 ;
        RECT 100.195 120.715 100.365 120.905 ;
        RECT 103.875 120.695 104.045 120.885 ;
        RECT 105.715 120.715 105.885 120.905 ;
        RECT 107.550 120.745 107.670 120.855 ;
        RECT 108.935 120.695 109.105 120.905 ;
        RECT 35.195 119.885 36.565 120.695 ;
        RECT 36.575 119.885 42.085 120.695 ;
        RECT 42.095 119.885 47.605 120.695 ;
        RECT 47.615 119.885 53.125 120.695 ;
        RECT 53.135 119.885 58.645 120.695 ;
        RECT 58.655 119.885 60.485 120.695 ;
        RECT 60.965 119.825 61.395 120.610 ;
        RECT 61.415 119.885 66.925 120.695 ;
        RECT 66.935 119.885 72.445 120.695 ;
        RECT 72.455 119.885 77.965 120.695 ;
        RECT 77.975 119.885 83.485 120.695 ;
        RECT 83.495 119.885 86.245 120.695 ;
        RECT 86.725 119.825 87.155 120.610 ;
        RECT 87.175 119.885 92.685 120.695 ;
        RECT 92.695 119.885 98.205 120.695 ;
        RECT 98.215 119.885 103.725 120.695 ;
        RECT 103.735 119.885 107.405 120.695 ;
        RECT 107.875 119.885 109.245 120.695 ;
      LAYER nwell ;
        RECT 35.000 116.665 109.440 119.495 ;
      LAYER pwell ;
        RECT 35.195 115.465 36.565 116.275 ;
        RECT 36.575 115.465 42.085 116.275 ;
        RECT 42.095 115.465 47.605 116.275 ;
        RECT 48.085 115.550 48.515 116.335 ;
        RECT 48.535 115.465 54.045 116.275 ;
        RECT 54.055 115.465 59.565 116.275 ;
        RECT 59.575 115.465 65.085 116.275 ;
        RECT 65.095 115.465 70.605 116.275 ;
        RECT 70.615 115.465 73.365 116.275 ;
        RECT 73.845 115.550 74.275 116.335 ;
        RECT 74.295 115.465 79.805 116.275 ;
        RECT 79.815 115.465 85.325 116.275 ;
        RECT 85.335 115.465 90.845 116.275 ;
        RECT 90.855 115.465 96.365 116.275 ;
        RECT 96.375 115.465 99.125 116.275 ;
        RECT 99.605 115.550 100.035 116.335 ;
        RECT 100.055 115.465 105.565 116.275 ;
        RECT 105.575 115.465 107.405 116.275 ;
        RECT 107.875 115.465 109.245 116.275 ;
        RECT 35.335 115.255 35.505 115.465 ;
        RECT 36.715 115.255 36.885 115.465 ;
        RECT 42.235 115.255 42.405 115.465 ;
        RECT 47.755 115.415 47.925 115.445 ;
        RECT 47.750 115.305 47.925 115.415 ;
        RECT 47.755 115.255 47.925 115.305 ;
        RECT 48.675 115.275 48.845 115.465 ;
        RECT 53.275 115.255 53.445 115.445 ;
        RECT 54.195 115.275 54.365 115.465 ;
        RECT 58.795 115.255 58.965 115.445 ;
        RECT 59.715 115.275 59.885 115.465 ;
        RECT 60.630 115.305 60.750 115.415 ;
        RECT 61.555 115.255 61.725 115.445 ;
        RECT 65.235 115.275 65.405 115.465 ;
        RECT 67.075 115.255 67.245 115.445 ;
        RECT 70.755 115.275 70.925 115.465 ;
        RECT 72.595 115.255 72.765 115.445 ;
        RECT 73.510 115.305 73.630 115.415 ;
        RECT 74.435 115.275 74.605 115.465 ;
        RECT 78.115 115.255 78.285 115.445 ;
        RECT 79.955 115.275 80.125 115.465 ;
        RECT 83.635 115.255 83.805 115.445 ;
        RECT 85.475 115.275 85.645 115.465 ;
        RECT 86.390 115.305 86.510 115.415 ;
        RECT 87.315 115.255 87.485 115.445 ;
        RECT 90.995 115.275 91.165 115.465 ;
        RECT 92.835 115.255 93.005 115.445 ;
        RECT 96.515 115.275 96.685 115.465 ;
        RECT 98.355 115.255 98.525 115.445 ;
        RECT 99.270 115.305 99.390 115.415 ;
        RECT 100.195 115.275 100.365 115.465 ;
        RECT 103.875 115.255 104.045 115.445 ;
        RECT 105.715 115.275 105.885 115.465 ;
        RECT 107.550 115.305 107.670 115.415 ;
        RECT 108.935 115.255 109.105 115.465 ;
        RECT 35.195 114.445 36.565 115.255 ;
        RECT 36.575 114.445 42.085 115.255 ;
        RECT 42.095 114.445 47.605 115.255 ;
        RECT 47.615 114.445 53.125 115.255 ;
        RECT 53.135 114.445 58.645 115.255 ;
        RECT 58.655 114.445 60.485 115.255 ;
        RECT 60.965 114.385 61.395 115.170 ;
        RECT 61.415 114.445 66.925 115.255 ;
        RECT 66.935 114.445 72.445 115.255 ;
        RECT 72.455 114.445 77.965 115.255 ;
        RECT 77.975 114.445 83.485 115.255 ;
        RECT 83.495 114.445 86.245 115.255 ;
        RECT 86.725 114.385 87.155 115.170 ;
        RECT 87.175 114.445 92.685 115.255 ;
        RECT 92.695 114.445 98.205 115.255 ;
        RECT 98.215 114.445 103.725 115.255 ;
        RECT 103.735 114.445 107.405 115.255 ;
        RECT 107.875 114.445 109.245 115.255 ;
      LAYER nwell ;
        RECT 35.000 111.225 109.440 114.055 ;
      LAYER pwell ;
        RECT 35.195 110.025 36.565 110.835 ;
        RECT 36.575 110.025 42.085 110.835 ;
        RECT 42.095 110.025 47.605 110.835 ;
        RECT 48.085 110.110 48.515 110.895 ;
        RECT 48.535 110.025 54.045 110.835 ;
        RECT 54.055 110.025 59.565 110.835 ;
        RECT 59.575 110.025 65.085 110.835 ;
        RECT 65.095 110.025 70.605 110.835 ;
        RECT 70.615 110.025 73.365 110.835 ;
        RECT 73.845 110.110 74.275 110.895 ;
        RECT 74.295 110.025 79.805 110.835 ;
        RECT 79.815 110.025 85.325 110.835 ;
        RECT 85.335 110.025 90.845 110.835 ;
        RECT 90.855 110.025 96.365 110.835 ;
        RECT 96.375 110.025 99.125 110.835 ;
        RECT 99.605 110.110 100.035 110.895 ;
        RECT 100.055 110.025 105.565 110.835 ;
        RECT 105.575 110.025 107.405 110.835 ;
        RECT 107.875 110.025 109.245 110.835 ;
        RECT 35.335 109.815 35.505 110.025 ;
        RECT 36.715 109.815 36.885 110.025 ;
        RECT 42.235 109.815 42.405 110.025 ;
        RECT 47.755 109.975 47.925 110.005 ;
        RECT 47.750 109.865 47.925 109.975 ;
        RECT 47.755 109.815 47.925 109.865 ;
        RECT 48.675 109.835 48.845 110.025 ;
        RECT 53.275 109.815 53.445 110.005 ;
        RECT 54.195 109.835 54.365 110.025 ;
        RECT 58.795 109.815 58.965 110.005 ;
        RECT 59.715 109.835 59.885 110.025 ;
        RECT 60.630 109.865 60.750 109.975 ;
        RECT 61.555 109.815 61.725 110.005 ;
        RECT 65.235 109.835 65.405 110.025 ;
        RECT 67.075 109.815 67.245 110.005 ;
        RECT 70.755 109.835 70.925 110.025 ;
        RECT 72.595 109.815 72.765 110.005 ;
        RECT 73.510 109.865 73.630 109.975 ;
        RECT 74.435 109.835 74.605 110.025 ;
        RECT 78.115 109.815 78.285 110.005 ;
        RECT 79.955 109.835 80.125 110.025 ;
        RECT 83.635 109.815 83.805 110.005 ;
        RECT 85.475 109.835 85.645 110.025 ;
        RECT 86.390 109.865 86.510 109.975 ;
        RECT 87.315 109.815 87.485 110.005 ;
        RECT 90.995 109.835 91.165 110.025 ;
        RECT 92.835 109.815 93.005 110.005 ;
        RECT 96.515 109.835 96.685 110.025 ;
        RECT 98.355 109.815 98.525 110.005 ;
        RECT 99.270 109.865 99.390 109.975 ;
        RECT 100.195 109.835 100.365 110.025 ;
        RECT 103.875 109.815 104.045 110.005 ;
        RECT 105.715 109.835 105.885 110.025 ;
        RECT 107.550 109.865 107.670 109.975 ;
        RECT 108.935 109.815 109.105 110.025 ;
        RECT 35.195 109.005 36.565 109.815 ;
        RECT 36.575 109.005 42.085 109.815 ;
        RECT 42.095 109.005 47.605 109.815 ;
        RECT 47.615 109.005 53.125 109.815 ;
        RECT 53.135 109.005 58.645 109.815 ;
        RECT 58.655 109.005 60.485 109.815 ;
        RECT 60.965 108.945 61.395 109.730 ;
        RECT 61.415 109.005 66.925 109.815 ;
        RECT 66.935 109.005 72.445 109.815 ;
        RECT 72.455 109.005 77.965 109.815 ;
        RECT 77.975 109.005 83.485 109.815 ;
        RECT 83.495 109.005 86.245 109.815 ;
        RECT 86.725 108.945 87.155 109.730 ;
        RECT 87.175 109.005 92.685 109.815 ;
        RECT 92.695 109.005 98.205 109.815 ;
        RECT 98.215 109.005 103.725 109.815 ;
        RECT 103.735 109.005 107.405 109.815 ;
        RECT 107.875 109.005 109.245 109.815 ;
      LAYER nwell ;
        RECT 35.000 105.785 109.440 108.615 ;
      LAYER pwell ;
        RECT 35.195 104.585 36.565 105.395 ;
        RECT 36.575 104.585 42.085 105.395 ;
        RECT 42.095 104.585 47.605 105.395 ;
        RECT 48.085 104.670 48.515 105.455 ;
        RECT 48.535 104.585 54.045 105.395 ;
        RECT 54.055 104.585 59.565 105.395 ;
        RECT 59.575 104.585 65.085 105.395 ;
        RECT 65.095 104.585 70.605 105.395 ;
        RECT 70.615 104.585 73.365 105.395 ;
        RECT 73.845 104.670 74.275 105.455 ;
        RECT 74.295 104.585 79.805 105.395 ;
        RECT 79.815 104.585 85.325 105.395 ;
        RECT 85.335 104.585 90.845 105.395 ;
        RECT 90.855 104.585 96.365 105.395 ;
        RECT 96.375 104.585 99.125 105.395 ;
        RECT 99.605 104.670 100.035 105.455 ;
        RECT 100.055 104.585 105.565 105.395 ;
        RECT 105.575 104.585 107.405 105.395 ;
        RECT 107.875 104.585 109.245 105.395 ;
        RECT 35.335 104.375 35.505 104.585 ;
        RECT 36.715 104.375 36.885 104.585 ;
        RECT 42.235 104.375 42.405 104.585 ;
        RECT 47.755 104.535 47.925 104.565 ;
        RECT 47.750 104.425 47.925 104.535 ;
        RECT 47.755 104.375 47.925 104.425 ;
        RECT 48.675 104.395 48.845 104.585 ;
        RECT 53.275 104.375 53.445 104.565 ;
        RECT 54.195 104.395 54.365 104.585 ;
        RECT 58.795 104.375 58.965 104.565 ;
        RECT 59.715 104.395 59.885 104.585 ;
        RECT 60.630 104.425 60.750 104.535 ;
        RECT 61.555 104.375 61.725 104.565 ;
        RECT 65.235 104.395 65.405 104.585 ;
        RECT 67.075 104.375 67.245 104.565 ;
        RECT 70.755 104.395 70.925 104.585 ;
        RECT 72.595 104.375 72.765 104.565 ;
        RECT 73.510 104.425 73.630 104.535 ;
        RECT 74.435 104.395 74.605 104.585 ;
        RECT 78.115 104.375 78.285 104.565 ;
        RECT 79.955 104.395 80.125 104.585 ;
        RECT 83.635 104.375 83.805 104.565 ;
        RECT 85.475 104.395 85.645 104.585 ;
        RECT 86.390 104.425 86.510 104.535 ;
        RECT 87.315 104.375 87.485 104.565 ;
        RECT 90.995 104.395 91.165 104.585 ;
        RECT 92.835 104.375 93.005 104.565 ;
        RECT 96.515 104.395 96.685 104.585 ;
        RECT 98.355 104.375 98.525 104.565 ;
        RECT 99.270 104.425 99.390 104.535 ;
        RECT 100.195 104.395 100.365 104.585 ;
        RECT 103.875 104.375 104.045 104.565 ;
        RECT 105.715 104.395 105.885 104.585 ;
        RECT 107.550 104.425 107.670 104.535 ;
        RECT 108.935 104.375 109.105 104.585 ;
        RECT 35.195 103.565 36.565 104.375 ;
        RECT 36.575 103.565 42.085 104.375 ;
        RECT 42.095 103.565 47.605 104.375 ;
        RECT 47.615 103.565 53.125 104.375 ;
        RECT 53.135 103.565 58.645 104.375 ;
        RECT 58.655 103.565 60.485 104.375 ;
        RECT 60.965 103.505 61.395 104.290 ;
        RECT 61.415 103.565 66.925 104.375 ;
        RECT 66.935 103.565 72.445 104.375 ;
        RECT 72.455 103.565 77.965 104.375 ;
        RECT 77.975 103.565 83.485 104.375 ;
        RECT 83.495 103.565 86.245 104.375 ;
        RECT 86.725 103.505 87.155 104.290 ;
        RECT 87.175 103.565 92.685 104.375 ;
        RECT 92.695 103.565 98.205 104.375 ;
        RECT 98.215 103.565 103.725 104.375 ;
        RECT 103.735 103.565 107.405 104.375 ;
        RECT 107.875 103.565 109.245 104.375 ;
      LAYER nwell ;
        RECT 35.000 100.345 109.440 103.175 ;
      LAYER pwell ;
        RECT 35.195 99.145 36.565 99.955 ;
        RECT 36.575 99.145 42.085 99.955 ;
        RECT 42.095 99.145 47.605 99.955 ;
        RECT 48.085 99.230 48.515 100.015 ;
        RECT 48.535 99.145 54.045 99.955 ;
        RECT 54.055 99.145 59.565 99.955 ;
        RECT 59.575 99.145 65.085 99.955 ;
        RECT 65.095 99.145 70.605 99.955 ;
        RECT 70.615 99.145 73.365 99.955 ;
        RECT 73.845 99.230 74.275 100.015 ;
        RECT 74.295 99.145 79.805 99.955 ;
        RECT 79.815 99.145 85.325 99.955 ;
        RECT 85.335 99.145 90.845 99.955 ;
        RECT 90.855 99.145 96.365 99.955 ;
        RECT 96.375 99.145 99.125 99.955 ;
        RECT 99.605 99.230 100.035 100.015 ;
        RECT 100.055 99.145 105.565 99.955 ;
        RECT 105.575 99.145 107.405 99.955 ;
        RECT 107.875 99.145 109.245 99.955 ;
        RECT 35.335 98.935 35.505 99.145 ;
        RECT 36.715 98.935 36.885 99.145 ;
        RECT 42.235 98.935 42.405 99.145 ;
        RECT 47.755 99.095 47.925 99.125 ;
        RECT 47.750 98.985 47.925 99.095 ;
        RECT 47.755 98.935 47.925 98.985 ;
        RECT 48.675 98.955 48.845 99.145 ;
        RECT 53.275 98.935 53.445 99.125 ;
        RECT 54.195 98.955 54.365 99.145 ;
        RECT 58.795 98.935 58.965 99.125 ;
        RECT 59.715 98.955 59.885 99.145 ;
        RECT 60.630 98.985 60.750 99.095 ;
        RECT 61.555 98.935 61.725 99.125 ;
        RECT 65.235 98.955 65.405 99.145 ;
        RECT 67.075 98.935 67.245 99.125 ;
        RECT 70.755 98.955 70.925 99.145 ;
        RECT 72.595 98.935 72.765 99.125 ;
        RECT 73.510 98.985 73.630 99.095 ;
        RECT 74.435 98.955 74.605 99.145 ;
        RECT 78.115 98.935 78.285 99.125 ;
        RECT 79.955 98.955 80.125 99.145 ;
        RECT 83.635 98.935 83.805 99.125 ;
        RECT 85.475 98.955 85.645 99.145 ;
        RECT 86.390 98.985 86.510 99.095 ;
        RECT 87.315 98.935 87.485 99.125 ;
        RECT 90.995 98.955 91.165 99.145 ;
        RECT 92.835 98.935 93.005 99.125 ;
        RECT 96.515 98.955 96.685 99.145 ;
        RECT 98.355 98.935 98.525 99.125 ;
        RECT 99.270 98.985 99.390 99.095 ;
        RECT 100.195 98.955 100.365 99.145 ;
        RECT 103.875 98.935 104.045 99.125 ;
        RECT 105.715 98.955 105.885 99.145 ;
        RECT 107.550 98.985 107.670 99.095 ;
        RECT 108.935 98.935 109.105 99.145 ;
        RECT 35.195 98.125 36.565 98.935 ;
        RECT 36.575 98.125 42.085 98.935 ;
        RECT 42.095 98.125 47.605 98.935 ;
        RECT 47.615 98.125 53.125 98.935 ;
        RECT 53.135 98.125 58.645 98.935 ;
        RECT 58.655 98.125 60.485 98.935 ;
        RECT 60.965 98.065 61.395 98.850 ;
        RECT 61.415 98.125 66.925 98.935 ;
        RECT 66.935 98.125 72.445 98.935 ;
        RECT 72.455 98.125 77.965 98.935 ;
        RECT 77.975 98.125 83.485 98.935 ;
        RECT 83.495 98.125 86.245 98.935 ;
        RECT 86.725 98.065 87.155 98.850 ;
        RECT 87.175 98.125 92.685 98.935 ;
        RECT 92.695 98.125 98.205 98.935 ;
        RECT 98.215 98.125 103.725 98.935 ;
        RECT 103.735 98.125 107.405 98.935 ;
        RECT 107.875 98.125 109.245 98.935 ;
      LAYER nwell ;
        RECT 35.000 94.905 109.440 97.735 ;
      LAYER pwell ;
        RECT 35.195 93.705 36.565 94.515 ;
        RECT 36.575 93.705 42.085 94.515 ;
        RECT 42.095 93.705 47.605 94.515 ;
        RECT 48.085 93.790 48.515 94.575 ;
        RECT 48.535 93.705 54.045 94.515 ;
        RECT 54.055 93.705 59.565 94.515 ;
        RECT 59.575 93.705 65.085 94.515 ;
        RECT 65.095 93.705 70.605 94.515 ;
        RECT 70.615 93.705 73.365 94.515 ;
        RECT 73.845 93.790 74.275 94.575 ;
        RECT 74.295 93.705 79.805 94.515 ;
        RECT 79.815 93.705 85.325 94.515 ;
        RECT 85.335 93.705 90.845 94.515 ;
        RECT 90.855 93.705 96.365 94.515 ;
        RECT 96.375 93.705 99.125 94.515 ;
        RECT 99.605 93.790 100.035 94.575 ;
        RECT 100.055 93.705 105.565 94.515 ;
        RECT 105.575 93.705 107.405 94.515 ;
        RECT 107.875 93.705 109.245 94.515 ;
        RECT 35.335 93.495 35.505 93.705 ;
        RECT 36.715 93.495 36.885 93.705 ;
        RECT 42.235 93.495 42.405 93.705 ;
        RECT 47.755 93.655 47.925 93.685 ;
        RECT 47.750 93.545 47.925 93.655 ;
        RECT 47.755 93.495 47.925 93.545 ;
        RECT 48.675 93.515 48.845 93.705 ;
        RECT 53.275 93.495 53.445 93.685 ;
        RECT 54.195 93.515 54.365 93.705 ;
        RECT 58.795 93.495 58.965 93.685 ;
        RECT 59.715 93.515 59.885 93.705 ;
        RECT 60.630 93.545 60.750 93.655 ;
        RECT 61.555 93.495 61.725 93.685 ;
        RECT 65.235 93.515 65.405 93.705 ;
        RECT 67.075 93.495 67.245 93.685 ;
        RECT 70.755 93.515 70.925 93.705 ;
        RECT 72.595 93.495 72.765 93.685 ;
        RECT 73.510 93.545 73.630 93.655 ;
        RECT 74.435 93.515 74.605 93.705 ;
        RECT 78.115 93.495 78.285 93.685 ;
        RECT 79.955 93.515 80.125 93.705 ;
        RECT 83.635 93.495 83.805 93.685 ;
        RECT 85.475 93.515 85.645 93.705 ;
        RECT 86.390 93.545 86.510 93.655 ;
        RECT 87.315 93.495 87.485 93.685 ;
        RECT 90.995 93.515 91.165 93.705 ;
        RECT 92.835 93.495 93.005 93.685 ;
        RECT 96.515 93.515 96.685 93.705 ;
        RECT 98.355 93.495 98.525 93.685 ;
        RECT 99.270 93.545 99.390 93.655 ;
        RECT 100.195 93.515 100.365 93.705 ;
        RECT 103.875 93.495 104.045 93.685 ;
        RECT 105.715 93.515 105.885 93.705 ;
        RECT 107.550 93.545 107.670 93.655 ;
        RECT 108.935 93.495 109.105 93.705 ;
        RECT 35.195 92.685 36.565 93.495 ;
        RECT 36.575 92.685 42.085 93.495 ;
        RECT 42.095 92.685 47.605 93.495 ;
        RECT 47.615 92.685 53.125 93.495 ;
        RECT 53.135 92.685 58.645 93.495 ;
        RECT 58.655 92.685 60.485 93.495 ;
        RECT 60.965 92.625 61.395 93.410 ;
        RECT 61.415 92.685 66.925 93.495 ;
        RECT 66.935 92.685 72.445 93.495 ;
        RECT 72.455 92.685 77.965 93.495 ;
        RECT 77.975 92.685 83.485 93.495 ;
        RECT 83.495 92.685 86.245 93.495 ;
        RECT 86.725 92.625 87.155 93.410 ;
        RECT 87.175 92.685 92.685 93.495 ;
        RECT 92.695 92.685 98.205 93.495 ;
        RECT 98.215 92.685 103.725 93.495 ;
        RECT 103.735 92.685 107.405 93.495 ;
        RECT 107.875 92.685 109.245 93.495 ;
      LAYER nwell ;
        RECT 35.000 89.465 109.440 92.295 ;
      LAYER pwell ;
        RECT 35.195 88.265 36.565 89.075 ;
        RECT 36.575 88.265 42.085 89.075 ;
        RECT 42.095 88.265 47.605 89.075 ;
        RECT 48.085 88.350 48.515 89.135 ;
        RECT 48.535 88.265 54.045 89.075 ;
        RECT 54.055 88.265 59.565 89.075 ;
        RECT 59.575 88.265 65.085 89.075 ;
        RECT 65.095 88.265 70.605 89.075 ;
        RECT 70.615 88.265 73.365 89.075 ;
        RECT 73.845 88.350 74.275 89.135 ;
        RECT 74.295 88.265 79.805 89.075 ;
        RECT 79.815 88.265 85.325 89.075 ;
        RECT 85.335 88.265 90.845 89.075 ;
        RECT 90.855 88.265 96.365 89.075 ;
        RECT 96.375 88.265 99.125 89.075 ;
        RECT 99.605 88.350 100.035 89.135 ;
        RECT 100.055 88.265 105.565 89.075 ;
        RECT 105.575 88.265 107.405 89.075 ;
        RECT 107.875 88.265 109.245 89.075 ;
        RECT 35.335 88.055 35.505 88.265 ;
        RECT 36.715 88.055 36.885 88.265 ;
        RECT 42.235 88.055 42.405 88.265 ;
        RECT 47.755 88.215 47.925 88.245 ;
        RECT 47.750 88.105 47.925 88.215 ;
        RECT 47.755 88.055 47.925 88.105 ;
        RECT 48.675 88.075 48.845 88.265 ;
        RECT 53.275 88.055 53.445 88.245 ;
        RECT 54.195 88.075 54.365 88.265 ;
        RECT 58.795 88.055 58.965 88.245 ;
        RECT 59.715 88.075 59.885 88.265 ;
        RECT 60.630 88.105 60.750 88.215 ;
        RECT 61.555 88.055 61.725 88.245 ;
        RECT 65.235 88.075 65.405 88.265 ;
        RECT 67.075 88.055 67.245 88.245 ;
        RECT 70.755 88.075 70.925 88.265 ;
        RECT 72.595 88.055 72.765 88.245 ;
        RECT 73.510 88.105 73.630 88.215 ;
        RECT 74.435 88.075 74.605 88.265 ;
        RECT 78.115 88.055 78.285 88.245 ;
        RECT 79.955 88.075 80.125 88.265 ;
        RECT 83.635 88.055 83.805 88.245 ;
        RECT 85.475 88.075 85.645 88.265 ;
        RECT 86.390 88.105 86.510 88.215 ;
        RECT 87.315 88.055 87.485 88.245 ;
        RECT 90.995 88.075 91.165 88.265 ;
        RECT 92.835 88.055 93.005 88.245 ;
        RECT 96.515 88.075 96.685 88.265 ;
        RECT 98.355 88.055 98.525 88.245 ;
        RECT 99.270 88.105 99.390 88.215 ;
        RECT 100.195 88.075 100.365 88.265 ;
        RECT 103.875 88.055 104.045 88.245 ;
        RECT 105.715 88.075 105.885 88.265 ;
        RECT 107.550 88.105 107.670 88.215 ;
        RECT 108.935 88.055 109.105 88.265 ;
        RECT 35.195 87.245 36.565 88.055 ;
        RECT 36.575 87.245 42.085 88.055 ;
        RECT 42.095 87.245 47.605 88.055 ;
        RECT 47.615 87.245 53.125 88.055 ;
        RECT 53.135 87.245 58.645 88.055 ;
        RECT 58.655 87.245 60.485 88.055 ;
        RECT 60.965 87.185 61.395 87.970 ;
        RECT 61.415 87.245 66.925 88.055 ;
        RECT 66.935 87.245 72.445 88.055 ;
        RECT 72.455 87.245 77.965 88.055 ;
        RECT 77.975 87.245 83.485 88.055 ;
        RECT 83.495 87.245 86.245 88.055 ;
        RECT 86.725 87.185 87.155 87.970 ;
        RECT 87.175 87.245 92.685 88.055 ;
        RECT 92.695 87.245 98.205 88.055 ;
        RECT 98.215 87.245 103.725 88.055 ;
        RECT 103.735 87.245 107.405 88.055 ;
        RECT 107.875 87.245 109.245 88.055 ;
      LAYER nwell ;
        RECT 35.000 84.025 109.440 86.855 ;
      LAYER pwell ;
        RECT 35.195 82.825 36.565 83.635 ;
        RECT 36.575 82.825 42.085 83.635 ;
        RECT 42.095 82.825 47.605 83.635 ;
        RECT 48.085 82.910 48.515 83.695 ;
        RECT 48.535 82.825 54.045 83.635 ;
        RECT 54.055 82.825 59.565 83.635 ;
        RECT 59.575 82.825 60.945 83.635 ;
        RECT 60.965 82.910 61.395 83.695 ;
        RECT 61.415 82.825 66.925 83.635 ;
        RECT 66.935 82.825 72.445 83.635 ;
        RECT 72.455 82.825 73.825 83.635 ;
        RECT 73.845 82.910 74.275 83.695 ;
        RECT 74.295 82.825 76.125 83.505 ;
        RECT 76.135 82.825 81.645 83.635 ;
        RECT 81.655 82.825 85.325 83.635 ;
        RECT 85.335 82.825 86.705 83.635 ;
        RECT 86.725 82.910 87.155 83.695 ;
        RECT 87.175 82.825 92.685 83.635 ;
        RECT 92.695 82.825 98.205 83.635 ;
        RECT 98.215 82.825 99.585 83.635 ;
        RECT 99.605 82.910 100.035 83.695 ;
        RECT 100.055 82.825 105.565 83.635 ;
        RECT 105.575 82.825 107.405 83.635 ;
        RECT 107.875 82.825 109.245 83.635 ;
        RECT 35.335 82.635 35.505 82.825 ;
        RECT 36.715 82.635 36.885 82.825 ;
        RECT 42.235 82.635 42.405 82.825 ;
        RECT 47.750 82.665 47.870 82.775 ;
        RECT 48.675 82.635 48.845 82.825 ;
        RECT 54.195 82.635 54.365 82.825 ;
        RECT 59.715 82.635 59.885 82.825 ;
        RECT 61.555 82.635 61.725 82.825 ;
        RECT 67.075 82.635 67.245 82.825 ;
        RECT 72.595 82.635 72.765 82.825 ;
        RECT 74.435 82.635 74.605 82.825 ;
        RECT 76.275 82.635 76.445 82.825 ;
        RECT 81.795 82.635 81.965 82.825 ;
        RECT 85.475 82.635 85.645 82.825 ;
        RECT 87.315 82.635 87.485 82.825 ;
        RECT 92.835 82.635 93.005 82.825 ;
        RECT 98.355 82.635 98.525 82.825 ;
        RECT 100.195 82.635 100.365 82.825 ;
        RECT 105.715 82.635 105.885 82.825 ;
        RECT 107.550 82.665 107.670 82.775 ;
        RECT 108.935 82.635 109.105 82.825 ;
      LAYER nwell ;
        RECT 110.050 77.920 136.970 77.930 ;
        RECT 21.800 69.100 37.850 73.650 ;
        RECT 40.000 65.400 104.800 72.000 ;
        RECT 40.000 41.850 96.700 65.400 ;
        RECT 106.350 59.310 136.970 77.920 ;
        RECT 106.350 59.300 111.010 59.310 ;
      LAYER pwell ;
        RECT 110.200 58.720 136.820 58.730 ;
        RECT 106.500 49.460 136.820 58.720 ;
        RECT 106.500 49.450 110.860 49.460 ;
        RECT 105.020 35.000 137.790 47.820 ;
      LAYER nwell ;
        RECT 20.050 27.450 95.700 31.850 ;
        RECT 20.050 22.450 83.750 27.450 ;
      LAYER li1 ;
        RECT 35.190 156.075 109.250 156.245 ;
        RECT 35.275 154.985 36.485 156.075 ;
        RECT 35.275 154.275 35.795 154.815 ;
        RECT 35.965 154.445 36.485 154.985 ;
        RECT 37.655 155.145 37.835 155.905 ;
        RECT 38.015 155.315 38.345 156.075 ;
        RECT 37.655 154.975 38.330 155.145 ;
        RECT 38.515 155.000 38.785 155.905 ;
        RECT 38.955 155.640 44.300 156.075 ;
        RECT 38.160 154.830 38.330 154.975 ;
        RECT 37.595 154.425 37.935 154.795 ;
        RECT 38.160 154.500 38.435 154.830 ;
        RECT 35.275 153.525 36.485 154.275 ;
        RECT 38.160 154.245 38.330 154.500 ;
        RECT 37.665 154.075 38.330 154.245 ;
        RECT 38.605 154.200 38.785 155.000 ;
        RECT 37.665 153.695 37.835 154.075 ;
        RECT 38.015 153.525 38.345 153.905 ;
        RECT 38.525 153.695 38.785 154.200 ;
        RECT 40.540 154.070 40.880 154.900 ;
        RECT 42.360 154.390 42.710 155.640 ;
        RECT 44.475 154.985 47.985 156.075 ;
        RECT 44.475 154.295 46.125 154.815 ;
        RECT 46.295 154.465 47.985 154.985 ;
        RECT 48.155 154.910 48.445 156.075 ;
        RECT 48.615 155.640 53.960 156.075 ;
        RECT 54.135 155.640 59.480 156.075 ;
        RECT 38.955 153.525 44.300 154.070 ;
        RECT 44.475 153.525 47.985 154.295 ;
        RECT 48.155 153.525 48.445 154.250 ;
        RECT 50.200 154.070 50.540 154.900 ;
        RECT 52.020 154.390 52.370 155.640 ;
        RECT 55.720 154.070 56.060 154.900 ;
        RECT 57.540 154.390 57.890 155.640 ;
        RECT 59.655 154.985 60.865 156.075 ;
        RECT 59.655 154.275 60.175 154.815 ;
        RECT 60.345 154.445 60.865 154.985 ;
        RECT 61.035 154.910 61.325 156.075 ;
        RECT 61.495 155.640 66.840 156.075 ;
        RECT 67.015 155.640 72.360 156.075 ;
        RECT 48.615 153.525 53.960 154.070 ;
        RECT 54.135 153.525 59.480 154.070 ;
        RECT 59.655 153.525 60.865 154.275 ;
        RECT 61.035 153.525 61.325 154.250 ;
        RECT 63.080 154.070 63.420 154.900 ;
        RECT 64.900 154.390 65.250 155.640 ;
        RECT 68.600 154.070 68.940 154.900 ;
        RECT 70.420 154.390 70.770 155.640 ;
        RECT 72.535 154.985 73.745 156.075 ;
        RECT 72.535 154.275 73.055 154.815 ;
        RECT 73.225 154.445 73.745 154.985 ;
        RECT 73.915 154.910 74.205 156.075 ;
        RECT 74.875 154.935 75.105 156.075 ;
        RECT 75.275 154.925 75.605 155.905 ;
        RECT 75.775 154.935 75.985 156.075 ;
        RECT 76.215 155.640 81.560 156.075 ;
        RECT 74.855 154.515 75.185 154.765 ;
        RECT 61.495 153.525 66.840 154.070 ;
        RECT 67.015 153.525 72.360 154.070 ;
        RECT 72.535 153.525 73.745 154.275 ;
        RECT 73.915 153.525 74.205 154.250 ;
        RECT 74.875 153.525 75.105 154.345 ;
        RECT 75.355 154.325 75.605 154.925 ;
        RECT 75.275 153.695 75.605 154.325 ;
        RECT 75.775 153.525 75.985 154.345 ;
        RECT 77.800 154.070 78.140 154.900 ;
        RECT 79.620 154.390 79.970 155.640 ;
        RECT 81.735 154.985 85.245 156.075 ;
        RECT 85.415 154.985 86.625 156.075 ;
        RECT 81.735 154.295 83.385 154.815 ;
        RECT 83.555 154.465 85.245 154.985 ;
        RECT 76.215 153.525 81.560 154.070 ;
        RECT 81.735 153.525 85.245 154.295 ;
        RECT 85.415 154.275 85.935 154.815 ;
        RECT 86.105 154.445 86.625 154.985 ;
        RECT 86.795 154.910 87.085 156.075 ;
        RECT 87.255 155.640 92.600 156.075 ;
        RECT 92.775 155.640 98.120 156.075 ;
        RECT 85.415 153.525 86.625 154.275 ;
        RECT 86.795 153.525 87.085 154.250 ;
        RECT 88.840 154.070 89.180 154.900 ;
        RECT 90.660 154.390 91.010 155.640 ;
        RECT 94.360 154.070 94.700 154.900 ;
        RECT 96.180 154.390 96.530 155.640 ;
        RECT 98.295 154.985 99.505 156.075 ;
        RECT 98.295 154.275 98.815 154.815 ;
        RECT 98.985 154.445 99.505 154.985 ;
        RECT 99.675 154.910 99.965 156.075 ;
        RECT 100.135 155.640 105.480 156.075 ;
        RECT 87.255 153.525 92.600 154.070 ;
        RECT 92.775 153.525 98.120 154.070 ;
        RECT 98.295 153.525 99.505 154.275 ;
        RECT 99.675 153.525 99.965 154.250 ;
        RECT 101.720 154.070 102.060 154.900 ;
        RECT 103.540 154.390 103.890 155.640 ;
        RECT 105.655 154.985 107.325 156.075 ;
        RECT 105.655 154.295 106.405 154.815 ;
        RECT 106.575 154.465 107.325 154.985 ;
        RECT 107.955 154.985 109.165 156.075 ;
        RECT 107.955 154.445 108.475 154.985 ;
        RECT 100.135 153.525 105.480 154.070 ;
        RECT 105.655 153.525 107.325 154.295 ;
        RECT 108.645 154.275 109.165 154.815 ;
        RECT 107.955 153.525 109.165 154.275 ;
        RECT 35.190 153.355 109.250 153.525 ;
        RECT 35.275 152.605 36.485 153.355 ;
        RECT 36.655 152.810 42.000 153.355 ;
        RECT 42.175 152.810 47.520 153.355 ;
        RECT 47.695 152.810 53.040 153.355 ;
        RECT 35.275 152.065 35.795 152.605 ;
        RECT 35.965 151.895 36.485 152.435 ;
        RECT 38.240 151.980 38.580 152.810 ;
        RECT 35.275 150.805 36.485 151.895 ;
        RECT 40.060 151.240 40.410 152.490 ;
        RECT 43.760 151.980 44.100 152.810 ;
        RECT 45.580 151.240 45.930 152.490 ;
        RECT 49.280 151.980 49.620 152.810 ;
        RECT 53.215 152.585 54.885 153.355 ;
        RECT 55.605 152.705 55.775 153.185 ;
        RECT 55.955 152.875 56.195 153.355 ;
        RECT 56.445 152.705 56.615 153.185 ;
        RECT 56.785 152.875 57.115 153.355 ;
        RECT 57.285 152.705 57.455 153.185 ;
        RECT 51.100 151.240 51.450 152.490 ;
        RECT 53.215 152.065 53.965 152.585 ;
        RECT 55.605 152.535 56.240 152.705 ;
        RECT 56.445 152.535 57.455 152.705 ;
        RECT 57.625 152.555 57.955 153.355 ;
        RECT 58.335 152.535 58.545 153.355 ;
        RECT 58.715 152.555 59.045 153.185 ;
        RECT 54.135 151.895 54.885 152.415 ;
        RECT 56.070 152.365 56.240 152.535 ;
        RECT 56.955 152.505 57.455 152.535 ;
        RECT 55.520 152.125 55.900 152.365 ;
        RECT 56.070 152.195 56.570 152.365 ;
        RECT 56.070 151.955 56.240 152.195 ;
        RECT 56.960 151.995 57.455 152.505 ;
        RECT 36.655 150.805 42.000 151.240 ;
        RECT 42.175 150.805 47.520 151.240 ;
        RECT 47.695 150.805 53.040 151.240 ;
        RECT 53.215 150.805 54.885 151.895 ;
        RECT 55.525 151.785 56.240 151.955 ;
        RECT 56.445 151.825 57.455 151.995 ;
        RECT 58.715 151.955 58.965 152.555 ;
        RECT 59.215 152.535 59.445 153.355 ;
        RECT 59.655 152.605 60.865 153.355 ;
        RECT 61.035 152.630 61.325 153.355 ;
        RECT 59.135 152.115 59.465 152.365 ;
        RECT 59.655 152.065 60.175 152.605 ;
        RECT 61.555 152.535 61.765 153.355 ;
        RECT 61.935 152.555 62.265 153.185 ;
        RECT 55.525 150.975 55.855 151.785 ;
        RECT 56.025 150.805 56.265 151.605 ;
        RECT 56.445 150.975 56.615 151.825 ;
        RECT 56.785 150.805 57.115 151.605 ;
        RECT 57.285 150.975 57.455 151.825 ;
        RECT 57.625 150.805 57.955 151.955 ;
        RECT 58.335 150.805 58.545 151.945 ;
        RECT 58.715 150.975 59.045 151.955 ;
        RECT 59.215 150.805 59.445 151.945 ;
        RECT 60.345 151.895 60.865 152.435 ;
        RECT 59.655 150.805 60.865 151.895 ;
        RECT 61.035 150.805 61.325 151.970 ;
        RECT 61.935 151.955 62.185 152.555 ;
        RECT 62.435 152.535 62.665 153.355 ;
        RECT 62.935 152.535 63.145 153.355 ;
        RECT 63.315 152.555 63.645 153.185 ;
        RECT 62.355 152.115 62.685 152.365 ;
        RECT 63.315 151.955 63.565 152.555 ;
        RECT 63.815 152.535 64.045 153.355 ;
        RECT 64.755 152.535 64.985 153.355 ;
        RECT 65.155 152.555 65.485 153.185 ;
        RECT 63.735 152.115 64.065 152.365 ;
        RECT 64.735 152.115 65.065 152.365 ;
        RECT 65.235 151.955 65.485 152.555 ;
        RECT 65.655 152.535 65.865 153.355 ;
        RECT 66.100 152.805 66.355 153.095 ;
        RECT 66.525 152.975 66.855 153.355 ;
        RECT 66.100 152.635 66.850 152.805 ;
        RECT 61.555 150.805 61.765 151.945 ;
        RECT 61.935 150.975 62.265 151.955 ;
        RECT 62.435 150.805 62.665 151.945 ;
        RECT 62.935 150.805 63.145 151.945 ;
        RECT 63.315 150.975 63.645 151.955 ;
        RECT 63.815 150.805 64.045 151.945 ;
        RECT 64.755 150.805 64.985 151.945 ;
        RECT 65.155 150.975 65.485 151.955 ;
        RECT 65.655 150.805 65.865 151.945 ;
        RECT 66.100 151.815 66.450 152.465 ;
        RECT 66.620 151.645 66.850 152.635 ;
        RECT 66.100 151.475 66.850 151.645 ;
        RECT 66.100 150.975 66.355 151.475 ;
        RECT 66.525 150.805 66.855 151.305 ;
        RECT 67.025 150.975 67.195 153.095 ;
        RECT 67.555 152.995 67.885 153.355 ;
        RECT 68.055 152.965 68.550 153.135 ;
        RECT 68.755 152.965 69.610 153.135 ;
        RECT 67.425 151.775 67.885 152.825 ;
        RECT 67.365 150.990 67.690 151.775 ;
        RECT 68.055 151.605 68.225 152.965 ;
        RECT 68.395 152.055 68.745 152.675 ;
        RECT 68.915 152.455 69.270 152.675 ;
        RECT 68.915 151.865 69.085 152.455 ;
        RECT 69.440 152.255 69.610 152.965 ;
        RECT 70.485 152.895 70.815 153.355 ;
        RECT 71.025 152.995 71.375 153.165 ;
        RECT 69.815 152.425 70.605 152.675 ;
        RECT 71.025 152.605 71.285 152.995 ;
        RECT 71.595 152.905 72.545 153.185 ;
        RECT 72.715 152.915 72.905 153.355 ;
        RECT 73.075 152.975 74.145 153.145 ;
        RECT 70.775 152.255 70.945 152.435 ;
        RECT 68.055 151.435 68.450 151.605 ;
        RECT 68.620 151.475 69.085 151.865 ;
        RECT 69.255 152.085 70.945 152.255 ;
        RECT 68.280 151.305 68.450 151.435 ;
        RECT 69.255 151.305 69.425 152.085 ;
        RECT 71.115 151.915 71.285 152.605 ;
        RECT 69.785 151.745 71.285 151.915 ;
        RECT 71.475 151.945 71.685 152.735 ;
        RECT 71.855 152.115 72.205 152.735 ;
        RECT 72.375 152.125 72.545 152.905 ;
        RECT 73.075 152.745 73.245 152.975 ;
        RECT 72.715 152.575 73.245 152.745 ;
        RECT 72.715 152.295 72.935 152.575 ;
        RECT 73.415 152.405 73.655 152.805 ;
        RECT 72.375 151.955 72.780 152.125 ;
        RECT 73.115 152.035 73.655 152.405 ;
        RECT 73.825 152.620 74.145 152.975 ;
        RECT 74.390 152.895 74.695 153.355 ;
        RECT 74.865 152.645 75.120 153.175 ;
        RECT 73.825 152.445 74.150 152.620 ;
        RECT 73.825 152.145 74.740 152.445 ;
        RECT 74.000 152.115 74.740 152.145 ;
        RECT 71.475 151.785 72.150 151.945 ;
        RECT 72.610 151.865 72.780 151.955 ;
        RECT 71.475 151.775 72.440 151.785 ;
        RECT 71.115 151.605 71.285 151.745 ;
        RECT 67.860 150.805 68.110 151.265 ;
        RECT 68.280 150.975 68.530 151.305 ;
        RECT 68.745 150.975 69.425 151.305 ;
        RECT 69.595 151.405 70.670 151.575 ;
        RECT 71.115 151.435 71.675 151.605 ;
        RECT 71.980 151.485 72.440 151.775 ;
        RECT 72.610 151.695 73.830 151.865 ;
        RECT 69.595 151.065 69.765 151.405 ;
        RECT 70.000 150.805 70.330 151.235 ;
        RECT 70.500 151.065 70.670 151.405 ;
        RECT 70.965 150.805 71.335 151.265 ;
        RECT 71.505 150.975 71.675 151.435 ;
        RECT 72.610 151.315 72.780 151.695 ;
        RECT 74.000 151.525 74.170 152.115 ;
        RECT 74.910 151.995 75.120 152.645 ;
        RECT 76.220 152.805 76.475 153.095 ;
        RECT 76.645 152.975 76.975 153.355 ;
        RECT 76.220 152.635 76.970 152.805 ;
        RECT 71.910 150.975 72.780 151.315 ;
        RECT 73.370 151.355 74.170 151.525 ;
        RECT 72.950 150.805 73.200 151.265 ;
        RECT 73.370 151.065 73.540 151.355 ;
        RECT 73.720 150.805 74.050 151.185 ;
        RECT 74.390 150.805 74.695 151.945 ;
        RECT 74.865 151.115 75.120 151.995 ;
        RECT 76.220 151.815 76.570 152.465 ;
        RECT 76.740 151.645 76.970 152.635 ;
        RECT 76.220 151.475 76.970 151.645 ;
        RECT 76.220 150.975 76.475 151.475 ;
        RECT 76.645 150.805 76.975 151.305 ;
        RECT 77.145 150.975 77.315 153.095 ;
        RECT 77.675 152.995 78.005 153.355 ;
        RECT 78.175 152.965 78.670 153.135 ;
        RECT 78.875 152.965 79.730 153.135 ;
        RECT 77.545 151.775 78.005 152.825 ;
        RECT 77.485 150.990 77.810 151.775 ;
        RECT 78.175 151.605 78.345 152.965 ;
        RECT 78.515 152.055 78.865 152.675 ;
        RECT 79.035 152.455 79.390 152.675 ;
        RECT 79.035 151.865 79.205 152.455 ;
        RECT 79.560 152.255 79.730 152.965 ;
        RECT 80.605 152.895 80.935 153.355 ;
        RECT 81.145 152.995 81.495 153.165 ;
        RECT 79.935 152.425 80.725 152.675 ;
        RECT 81.145 152.605 81.405 152.995 ;
        RECT 81.715 152.905 82.665 153.185 ;
        RECT 82.835 152.915 83.025 153.355 ;
        RECT 83.195 152.975 84.265 153.145 ;
        RECT 80.895 152.255 81.065 152.435 ;
        RECT 78.175 151.435 78.570 151.605 ;
        RECT 78.740 151.475 79.205 151.865 ;
        RECT 79.375 152.085 81.065 152.255 ;
        RECT 78.400 151.305 78.570 151.435 ;
        RECT 79.375 151.305 79.545 152.085 ;
        RECT 81.235 151.915 81.405 152.605 ;
        RECT 79.905 151.745 81.405 151.915 ;
        RECT 81.595 151.945 81.805 152.735 ;
        RECT 81.975 152.115 82.325 152.735 ;
        RECT 82.495 152.125 82.665 152.905 ;
        RECT 83.195 152.745 83.365 152.975 ;
        RECT 82.835 152.575 83.365 152.745 ;
        RECT 82.835 152.295 83.055 152.575 ;
        RECT 83.535 152.405 83.775 152.805 ;
        RECT 82.495 151.955 82.900 152.125 ;
        RECT 83.235 152.035 83.775 152.405 ;
        RECT 83.945 152.620 84.265 152.975 ;
        RECT 84.510 152.895 84.815 153.355 ;
        RECT 84.985 152.645 85.240 153.175 ;
        RECT 83.945 152.445 84.270 152.620 ;
        RECT 83.945 152.145 84.860 152.445 ;
        RECT 84.120 152.115 84.860 152.145 ;
        RECT 81.595 151.785 82.270 151.945 ;
        RECT 82.730 151.865 82.900 151.955 ;
        RECT 81.595 151.775 82.560 151.785 ;
        RECT 81.235 151.605 81.405 151.745 ;
        RECT 77.980 150.805 78.230 151.265 ;
        RECT 78.400 150.975 78.650 151.305 ;
        RECT 78.865 150.975 79.545 151.305 ;
        RECT 79.715 151.405 80.790 151.575 ;
        RECT 81.235 151.435 81.795 151.605 ;
        RECT 82.100 151.485 82.560 151.775 ;
        RECT 82.730 151.695 83.950 151.865 ;
        RECT 79.715 151.065 79.885 151.405 ;
        RECT 80.120 150.805 80.450 151.235 ;
        RECT 80.620 151.065 80.790 151.405 ;
        RECT 81.085 150.805 81.455 151.265 ;
        RECT 81.625 150.975 81.795 151.435 ;
        RECT 82.730 151.315 82.900 151.695 ;
        RECT 84.120 151.525 84.290 152.115 ;
        RECT 85.030 151.995 85.240 152.645 ;
        RECT 85.475 152.535 85.685 153.355 ;
        RECT 85.855 152.555 86.185 153.185 ;
        RECT 82.030 150.975 82.900 151.315 ;
        RECT 83.490 151.355 84.290 151.525 ;
        RECT 83.070 150.805 83.320 151.265 ;
        RECT 83.490 151.065 83.660 151.355 ;
        RECT 83.840 150.805 84.170 151.185 ;
        RECT 84.510 150.805 84.815 151.945 ;
        RECT 84.985 151.115 85.240 151.995 ;
        RECT 85.855 151.955 86.105 152.555 ;
        RECT 86.355 152.535 86.585 153.355 ;
        RECT 86.795 152.630 87.085 153.355 ;
        RECT 87.260 152.805 87.515 153.095 ;
        RECT 87.685 152.975 88.015 153.355 ;
        RECT 87.260 152.635 88.010 152.805 ;
        RECT 86.275 152.115 86.605 152.365 ;
        RECT 85.475 150.805 85.685 151.945 ;
        RECT 85.855 150.975 86.185 151.955 ;
        RECT 86.355 150.805 86.585 151.945 ;
        RECT 86.795 150.805 87.085 151.970 ;
        RECT 87.260 151.815 87.610 152.465 ;
        RECT 87.780 151.645 88.010 152.635 ;
        RECT 87.260 151.475 88.010 151.645 ;
        RECT 87.260 150.975 87.515 151.475 ;
        RECT 87.685 150.805 88.015 151.305 ;
        RECT 88.185 150.975 88.355 153.095 ;
        RECT 88.715 152.995 89.045 153.355 ;
        RECT 89.215 152.965 89.710 153.135 ;
        RECT 89.915 152.965 90.770 153.135 ;
        RECT 88.585 151.775 89.045 152.825 ;
        RECT 88.525 150.990 88.850 151.775 ;
        RECT 89.215 151.605 89.385 152.965 ;
        RECT 89.555 152.055 89.905 152.675 ;
        RECT 90.075 152.455 90.430 152.675 ;
        RECT 90.075 151.865 90.245 152.455 ;
        RECT 90.600 152.255 90.770 152.965 ;
        RECT 91.645 152.895 91.975 153.355 ;
        RECT 92.185 152.995 92.535 153.165 ;
        RECT 90.975 152.425 91.765 152.675 ;
        RECT 92.185 152.605 92.445 152.995 ;
        RECT 92.755 152.905 93.705 153.185 ;
        RECT 93.875 152.915 94.065 153.355 ;
        RECT 94.235 152.975 95.305 153.145 ;
        RECT 91.935 152.255 92.105 152.435 ;
        RECT 89.215 151.435 89.610 151.605 ;
        RECT 89.780 151.475 90.245 151.865 ;
        RECT 90.415 152.085 92.105 152.255 ;
        RECT 89.440 151.305 89.610 151.435 ;
        RECT 90.415 151.305 90.585 152.085 ;
        RECT 92.275 151.915 92.445 152.605 ;
        RECT 90.945 151.745 92.445 151.915 ;
        RECT 92.635 151.945 92.845 152.735 ;
        RECT 93.015 152.115 93.365 152.735 ;
        RECT 93.535 152.125 93.705 152.905 ;
        RECT 94.235 152.745 94.405 152.975 ;
        RECT 93.875 152.575 94.405 152.745 ;
        RECT 93.875 152.295 94.095 152.575 ;
        RECT 94.575 152.405 94.815 152.805 ;
        RECT 93.535 151.955 93.940 152.125 ;
        RECT 94.275 152.035 94.815 152.405 ;
        RECT 94.985 152.620 95.305 152.975 ;
        RECT 95.550 152.895 95.855 153.355 ;
        RECT 96.025 152.645 96.280 153.175 ;
        RECT 94.985 152.445 95.310 152.620 ;
        RECT 94.985 152.145 95.900 152.445 ;
        RECT 95.160 152.115 95.900 152.145 ;
        RECT 92.635 151.785 93.310 151.945 ;
        RECT 93.770 151.865 93.940 151.955 ;
        RECT 92.635 151.775 93.600 151.785 ;
        RECT 92.275 151.605 92.445 151.745 ;
        RECT 89.020 150.805 89.270 151.265 ;
        RECT 89.440 150.975 89.690 151.305 ;
        RECT 89.905 150.975 90.585 151.305 ;
        RECT 90.755 151.405 91.830 151.575 ;
        RECT 92.275 151.435 92.835 151.605 ;
        RECT 93.140 151.485 93.600 151.775 ;
        RECT 93.770 151.695 94.990 151.865 ;
        RECT 90.755 151.065 90.925 151.405 ;
        RECT 91.160 150.805 91.490 151.235 ;
        RECT 91.660 151.065 91.830 151.405 ;
        RECT 92.125 150.805 92.495 151.265 ;
        RECT 92.665 150.975 92.835 151.435 ;
        RECT 93.770 151.315 93.940 151.695 ;
        RECT 95.160 151.525 95.330 152.115 ;
        RECT 96.070 151.995 96.280 152.645 ;
        RECT 96.495 152.535 96.725 153.355 ;
        RECT 96.895 152.555 97.225 153.185 ;
        RECT 96.475 152.115 96.805 152.365 ;
        RECT 93.070 150.975 93.940 151.315 ;
        RECT 94.530 151.355 95.330 151.525 ;
        RECT 94.110 150.805 94.360 151.265 ;
        RECT 94.530 151.065 94.700 151.355 ;
        RECT 94.880 150.805 95.210 151.185 ;
        RECT 95.550 150.805 95.855 151.945 ;
        RECT 96.025 151.115 96.280 151.995 ;
        RECT 96.975 151.955 97.225 152.555 ;
        RECT 97.395 152.535 97.605 153.355 ;
        RECT 97.835 152.810 103.180 153.355 ;
        RECT 99.420 151.980 99.760 152.810 ;
        RECT 103.355 152.585 106.865 153.355 ;
        RECT 107.955 152.605 109.165 153.355 ;
        RECT 96.495 150.805 96.725 151.945 ;
        RECT 96.895 150.975 97.225 151.955 ;
        RECT 97.395 150.805 97.605 151.945 ;
        RECT 101.240 151.240 101.590 152.490 ;
        RECT 103.355 152.065 105.005 152.585 ;
        RECT 105.175 151.895 106.865 152.415 ;
        RECT 97.835 150.805 103.180 151.240 ;
        RECT 103.355 150.805 106.865 151.895 ;
        RECT 107.955 151.895 108.475 152.435 ;
        RECT 108.645 152.065 109.165 152.605 ;
        RECT 107.955 150.805 109.165 151.895 ;
        RECT 35.190 150.635 109.250 150.805 ;
        RECT 35.275 149.545 36.485 150.635 ;
        RECT 36.655 150.200 42.000 150.635 ;
        RECT 42.175 150.200 47.520 150.635 ;
        RECT 35.275 148.835 35.795 149.375 ;
        RECT 35.965 149.005 36.485 149.545 ;
        RECT 35.275 148.085 36.485 148.835 ;
        RECT 38.240 148.630 38.580 149.460 ;
        RECT 40.060 148.950 40.410 150.200 ;
        RECT 43.760 148.630 44.100 149.460 ;
        RECT 45.580 148.950 45.930 150.200 ;
        RECT 48.155 149.470 48.445 150.635 ;
        RECT 48.615 150.200 53.960 150.635 ;
        RECT 36.655 148.085 42.000 148.630 ;
        RECT 42.175 148.085 47.520 148.630 ;
        RECT 48.155 148.085 48.445 148.810 ;
        RECT 50.200 148.630 50.540 149.460 ;
        RECT 52.020 148.950 52.370 150.200 ;
        RECT 54.135 149.545 55.345 150.635 ;
        RECT 55.520 149.965 55.775 150.465 ;
        RECT 55.945 150.135 56.275 150.635 ;
        RECT 55.520 149.795 56.270 149.965 ;
        RECT 54.135 148.835 54.655 149.375 ;
        RECT 54.825 149.005 55.345 149.545 ;
        RECT 55.520 148.975 55.870 149.625 ;
        RECT 48.615 148.085 53.960 148.630 ;
        RECT 54.135 148.085 55.345 148.835 ;
        RECT 56.040 148.805 56.270 149.795 ;
        RECT 55.520 148.635 56.270 148.805 ;
        RECT 55.520 148.345 55.775 148.635 ;
        RECT 55.945 148.085 56.275 148.465 ;
        RECT 56.445 148.345 56.615 150.465 ;
        RECT 56.785 149.665 57.110 150.450 ;
        RECT 57.280 150.175 57.530 150.635 ;
        RECT 57.700 150.135 57.950 150.465 ;
        RECT 58.165 150.135 58.845 150.465 ;
        RECT 57.700 150.005 57.870 150.135 ;
        RECT 57.475 149.835 57.870 150.005 ;
        RECT 56.845 148.615 57.305 149.665 ;
        RECT 57.475 148.475 57.645 149.835 ;
        RECT 58.040 149.575 58.505 149.965 ;
        RECT 57.815 148.765 58.165 149.385 ;
        RECT 58.335 148.985 58.505 149.575 ;
        RECT 58.675 149.355 58.845 150.135 ;
        RECT 59.015 150.035 59.185 150.375 ;
        RECT 59.420 150.205 59.750 150.635 ;
        RECT 59.920 150.035 60.090 150.375 ;
        RECT 60.385 150.175 60.755 150.635 ;
        RECT 59.015 149.865 60.090 150.035 ;
        RECT 60.925 150.005 61.095 150.465 ;
        RECT 61.330 150.125 62.200 150.465 ;
        RECT 62.370 150.175 62.620 150.635 ;
        RECT 60.535 149.835 61.095 150.005 ;
        RECT 60.535 149.695 60.705 149.835 ;
        RECT 59.205 149.525 60.705 149.695 ;
        RECT 61.400 149.665 61.860 149.955 ;
        RECT 58.675 149.185 60.365 149.355 ;
        RECT 58.335 148.765 58.690 148.985 ;
        RECT 58.860 148.475 59.030 149.185 ;
        RECT 59.235 148.765 60.025 149.015 ;
        RECT 60.195 149.005 60.365 149.185 ;
        RECT 60.535 148.835 60.705 149.525 ;
        RECT 56.975 148.085 57.305 148.445 ;
        RECT 57.475 148.305 57.970 148.475 ;
        RECT 58.175 148.305 59.030 148.475 ;
        RECT 59.905 148.085 60.235 148.545 ;
        RECT 60.445 148.445 60.705 148.835 ;
        RECT 60.895 149.655 61.860 149.665 ;
        RECT 62.030 149.745 62.200 150.125 ;
        RECT 62.790 150.085 62.960 150.375 ;
        RECT 63.140 150.255 63.470 150.635 ;
        RECT 62.790 149.915 63.590 150.085 ;
        RECT 60.895 149.495 61.570 149.655 ;
        RECT 62.030 149.575 63.250 149.745 ;
        RECT 60.895 148.705 61.105 149.495 ;
        RECT 62.030 149.485 62.200 149.575 ;
        RECT 61.275 148.705 61.625 149.325 ;
        RECT 61.795 149.315 62.200 149.485 ;
        RECT 61.795 148.535 61.965 149.315 ;
        RECT 62.135 148.865 62.355 149.145 ;
        RECT 62.535 149.035 63.075 149.405 ;
        RECT 63.420 149.325 63.590 149.915 ;
        RECT 63.810 149.495 64.115 150.635 ;
        RECT 64.285 149.445 64.540 150.325 ;
        RECT 64.830 150.005 65.115 150.465 ;
        RECT 65.285 150.175 65.555 150.635 ;
        RECT 64.830 149.785 65.785 150.005 ;
        RECT 63.420 149.295 64.160 149.325 ;
        RECT 62.135 148.695 62.665 148.865 ;
        RECT 60.445 148.275 60.795 148.445 ;
        RECT 61.015 148.255 61.965 148.535 ;
        RECT 62.135 148.085 62.325 148.525 ;
        RECT 62.495 148.465 62.665 148.695 ;
        RECT 62.835 148.635 63.075 149.035 ;
        RECT 63.245 148.995 64.160 149.295 ;
        RECT 63.245 148.820 63.570 148.995 ;
        RECT 63.245 148.465 63.565 148.820 ;
        RECT 64.330 148.795 64.540 149.445 ;
        RECT 64.715 149.055 65.405 149.615 ;
        RECT 65.575 148.885 65.785 149.785 ;
        RECT 62.495 148.295 63.565 148.465 ;
        RECT 63.810 148.085 64.115 148.545 ;
        RECT 64.285 148.265 64.540 148.795 ;
        RECT 64.830 148.715 65.785 148.885 ;
        RECT 65.955 149.615 66.355 150.465 ;
        RECT 66.545 150.005 66.825 150.465 ;
        RECT 67.345 150.175 67.670 150.635 ;
        RECT 66.545 149.785 67.670 150.005 ;
        RECT 65.955 149.055 67.050 149.615 ;
        RECT 67.220 149.325 67.670 149.785 ;
        RECT 67.840 149.495 68.225 150.465 ;
        RECT 68.405 149.915 68.735 150.635 ;
        RECT 64.830 148.255 65.115 148.715 ;
        RECT 65.285 148.085 65.555 148.545 ;
        RECT 65.955 148.255 66.355 149.055 ;
        RECT 67.220 148.995 67.775 149.325 ;
        RECT 67.220 148.885 67.670 148.995 ;
        RECT 66.545 148.715 67.670 148.885 ;
        RECT 67.945 148.825 68.225 149.495 ;
        RECT 68.395 149.275 68.625 149.615 ;
        RECT 68.915 149.275 69.130 150.390 ;
        RECT 69.325 149.690 69.655 150.465 ;
        RECT 69.825 149.860 70.535 150.635 ;
        RECT 69.325 149.475 70.475 149.690 ;
        RECT 68.395 149.075 68.725 149.275 ;
        RECT 68.915 149.095 69.365 149.275 ;
        RECT 69.035 149.075 69.365 149.095 ;
        RECT 69.535 149.075 70.005 149.305 ;
        RECT 70.190 148.905 70.475 149.475 ;
        RECT 70.705 149.030 70.985 150.465 ;
        RECT 71.195 149.495 71.425 150.635 ;
        RECT 71.595 149.485 71.925 150.465 ;
        RECT 72.095 149.495 72.305 150.635 ;
        RECT 72.535 149.545 73.745 150.635 ;
        RECT 71.175 149.075 71.505 149.325 ;
        RECT 66.545 148.255 66.825 148.715 ;
        RECT 67.345 148.085 67.670 148.545 ;
        RECT 67.840 148.255 68.225 148.825 ;
        RECT 68.395 148.715 69.575 148.905 ;
        RECT 68.395 148.255 68.735 148.715 ;
        RECT 69.245 148.635 69.575 148.715 ;
        RECT 69.765 148.715 70.475 148.905 ;
        RECT 69.765 148.575 70.065 148.715 ;
        RECT 69.750 148.565 70.065 148.575 ;
        RECT 69.740 148.555 70.065 148.565 ;
        RECT 69.730 148.550 70.065 148.555 ;
        RECT 68.905 148.085 69.075 148.545 ;
        RECT 69.725 148.540 70.065 148.550 ;
        RECT 69.720 148.535 70.065 148.540 ;
        RECT 69.715 148.525 70.065 148.535 ;
        RECT 69.710 148.520 70.065 148.525 ;
        RECT 69.705 148.255 70.065 148.520 ;
        RECT 70.305 148.085 70.475 148.545 ;
        RECT 70.645 148.255 70.985 149.030 ;
        RECT 71.195 148.085 71.425 148.905 ;
        RECT 71.675 148.885 71.925 149.485 ;
        RECT 71.595 148.255 71.925 148.885 ;
        RECT 72.095 148.085 72.305 148.905 ;
        RECT 72.535 148.835 73.055 149.375 ;
        RECT 73.225 149.005 73.745 149.545 ;
        RECT 73.915 149.470 74.205 150.635 ;
        RECT 74.375 149.495 74.760 150.465 ;
        RECT 74.930 150.175 75.255 150.635 ;
        RECT 75.775 150.005 76.055 150.465 ;
        RECT 74.930 149.785 76.055 150.005 ;
        RECT 72.535 148.085 73.745 148.835 ;
        RECT 74.375 148.825 74.655 149.495 ;
        RECT 74.930 149.325 75.380 149.785 ;
        RECT 76.245 149.615 76.645 150.465 ;
        RECT 77.045 150.175 77.315 150.635 ;
        RECT 77.485 150.005 77.770 150.465 ;
        RECT 74.825 148.995 75.380 149.325 ;
        RECT 75.550 149.055 76.645 149.615 ;
        RECT 74.930 148.885 75.380 148.995 ;
        RECT 73.915 148.085 74.205 148.810 ;
        RECT 74.375 148.255 74.760 148.825 ;
        RECT 74.930 148.715 76.055 148.885 ;
        RECT 74.930 148.085 75.255 148.545 ;
        RECT 75.775 148.255 76.055 148.715 ;
        RECT 76.245 148.255 76.645 149.055 ;
        RECT 76.815 149.785 77.770 150.005 ;
        RECT 76.815 148.885 77.025 149.785 ;
        RECT 78.145 149.705 78.315 150.465 ;
        RECT 78.530 149.875 78.860 150.635 ;
        RECT 77.195 149.055 77.885 149.615 ;
        RECT 78.145 149.535 78.860 149.705 ;
        RECT 79.030 149.560 79.285 150.465 ;
        RECT 78.055 148.985 78.410 149.355 ;
        RECT 78.690 149.325 78.860 149.535 ;
        RECT 78.690 148.995 78.945 149.325 ;
        RECT 76.815 148.715 77.770 148.885 ;
        RECT 78.690 148.805 78.860 148.995 ;
        RECT 79.115 148.830 79.285 149.560 ;
        RECT 79.460 149.485 79.720 150.635 ;
        RECT 79.895 149.545 83.405 150.635 ;
        RECT 77.045 148.085 77.315 148.545 ;
        RECT 77.485 148.255 77.770 148.715 ;
        RECT 78.145 148.635 78.860 148.805 ;
        RECT 78.145 148.255 78.315 148.635 ;
        RECT 78.530 148.085 78.860 148.465 ;
        RECT 79.030 148.255 79.285 148.830 ;
        RECT 79.460 148.085 79.720 148.925 ;
        RECT 79.895 148.855 81.545 149.375 ;
        RECT 81.715 149.025 83.405 149.545 ;
        RECT 84.095 149.495 84.305 150.635 ;
        RECT 84.475 149.485 84.805 150.465 ;
        RECT 84.975 149.495 85.205 150.635 ;
        RECT 85.880 149.495 86.200 150.635 ;
        RECT 79.895 148.085 83.405 148.855 ;
        RECT 84.095 148.085 84.305 148.905 ;
        RECT 84.475 148.885 84.725 149.485 ;
        RECT 86.380 149.325 86.575 150.375 ;
        RECT 86.755 149.785 87.085 150.465 ;
        RECT 87.285 149.835 87.540 150.635 ;
        RECT 86.755 149.505 87.105 149.785 ;
        RECT 84.895 149.075 85.225 149.325 ;
        RECT 85.940 149.275 86.200 149.325 ;
        RECT 85.935 149.105 86.200 149.275 ;
        RECT 85.940 148.995 86.200 149.105 ;
        RECT 86.380 148.995 86.765 149.325 ;
        RECT 86.935 149.125 87.105 149.505 ;
        RECT 87.295 149.295 87.540 149.655 ;
        RECT 87.715 149.545 90.305 150.635 ;
        RECT 86.935 148.955 87.455 149.125 ;
        RECT 84.475 148.255 84.805 148.885 ;
        RECT 84.975 148.085 85.205 148.905 ;
        RECT 85.880 148.615 87.095 148.785 ;
        RECT 85.880 148.265 86.170 148.615 ;
        RECT 86.365 148.085 86.695 148.445 ;
        RECT 86.865 148.310 87.095 148.615 ;
        RECT 87.285 148.595 87.455 148.955 ;
        RECT 87.715 148.855 88.925 149.375 ;
        RECT 89.095 149.025 90.305 149.545 ;
        RECT 90.975 149.495 91.205 150.635 ;
        RECT 91.375 149.485 91.705 150.465 ;
        RECT 91.875 149.495 92.085 150.635 ;
        RECT 92.315 150.200 97.660 150.635 ;
        RECT 90.955 149.075 91.285 149.325 ;
        RECT 87.285 148.425 87.485 148.595 ;
        RECT 87.285 148.390 87.455 148.425 ;
        RECT 87.715 148.085 90.305 148.855 ;
        RECT 90.975 148.085 91.205 148.905 ;
        RECT 91.455 148.885 91.705 149.485 ;
        RECT 91.375 148.255 91.705 148.885 ;
        RECT 91.875 148.085 92.085 148.905 ;
        RECT 93.900 148.630 94.240 149.460 ;
        RECT 95.720 148.950 96.070 150.200 ;
        RECT 97.835 149.545 99.505 150.635 ;
        RECT 97.835 148.855 98.585 149.375 ;
        RECT 98.755 149.025 99.505 149.545 ;
        RECT 99.675 149.470 99.965 150.635 ;
        RECT 100.135 150.200 105.480 150.635 ;
        RECT 92.315 148.085 97.660 148.630 ;
        RECT 97.835 148.085 99.505 148.855 ;
        RECT 99.675 148.085 99.965 148.810 ;
        RECT 101.720 148.630 102.060 149.460 ;
        RECT 103.540 148.950 103.890 150.200 ;
        RECT 105.655 149.545 107.325 150.635 ;
        RECT 105.655 148.855 106.405 149.375 ;
        RECT 106.575 149.025 107.325 149.545 ;
        RECT 107.955 149.545 109.165 150.635 ;
        RECT 107.955 149.005 108.475 149.545 ;
        RECT 100.135 148.085 105.480 148.630 ;
        RECT 105.655 148.085 107.325 148.855 ;
        RECT 108.645 148.835 109.165 149.375 ;
        RECT 107.955 148.085 109.165 148.835 ;
        RECT 35.190 147.915 109.250 148.085 ;
        RECT 35.275 147.165 36.485 147.915 ;
        RECT 36.655 147.370 42.000 147.915 ;
        RECT 42.175 147.370 47.520 147.915 ;
        RECT 35.275 146.625 35.795 147.165 ;
        RECT 35.965 146.455 36.485 146.995 ;
        RECT 38.240 146.540 38.580 147.370 ;
        RECT 35.275 145.365 36.485 146.455 ;
        RECT 40.060 145.800 40.410 147.050 ;
        RECT 43.760 146.540 44.100 147.370 ;
        RECT 45.580 145.800 45.930 147.050 ;
        RECT 47.695 146.260 48.215 147.745 ;
        RECT 48.385 147.255 48.725 147.915 ;
        RECT 49.075 147.145 50.745 147.915 ;
        RECT 36.655 145.365 42.000 145.800 ;
        RECT 42.175 145.365 47.520 145.800 ;
        RECT 47.885 145.365 48.215 146.090 ;
        RECT 48.385 145.535 48.905 147.085 ;
        RECT 49.075 146.625 49.825 147.145 ;
        RECT 50.975 147.095 51.185 147.915 ;
        RECT 51.355 147.115 51.685 147.745 ;
        RECT 49.995 146.455 50.745 146.975 ;
        RECT 51.355 146.515 51.605 147.115 ;
        RECT 51.855 147.095 52.085 147.915 ;
        RECT 52.295 147.145 55.805 147.915 ;
        RECT 56.435 147.305 56.775 147.720 ;
        RECT 56.945 147.475 57.115 147.915 ;
        RECT 57.305 147.525 58.565 147.705 ;
        RECT 57.305 147.305 57.635 147.525 ;
        RECT 56.435 147.175 57.635 147.305 ;
        RECT 57.805 147.175 58.155 147.355 ;
        RECT 51.775 146.675 52.105 146.925 ;
        RECT 52.295 146.625 53.945 147.145 ;
        RECT 56.435 147.135 57.465 147.175 ;
        RECT 49.075 145.365 50.745 146.455 ;
        RECT 50.975 145.365 51.185 146.505 ;
        RECT 51.355 145.535 51.685 146.515 ;
        RECT 51.855 145.365 52.085 146.505 ;
        RECT 54.115 146.455 55.805 146.975 ;
        RECT 56.435 146.725 56.895 146.925 ;
        RECT 57.065 146.755 57.430 146.925 ;
        RECT 57.065 146.555 57.245 146.755 ;
        RECT 57.645 146.585 57.815 147.005 ;
        RECT 52.295 145.365 55.805 146.455 ;
        RECT 56.435 145.365 56.755 146.545 ;
        RECT 56.925 146.385 57.245 146.555 ;
        RECT 56.925 145.595 57.125 146.385 ;
        RECT 57.415 146.335 57.815 146.585 ;
        RECT 57.985 146.165 58.155 147.175 ;
        RECT 57.315 145.955 58.155 146.165 ;
        RECT 58.325 146.010 58.565 147.335 ;
        RECT 58.740 147.240 59.015 147.585 ;
        RECT 59.205 147.515 59.585 147.915 ;
        RECT 59.755 147.345 59.925 147.695 ;
        RECT 60.095 147.515 60.425 147.915 ;
        RECT 60.595 147.345 60.850 147.695 ;
        RECT 58.740 146.505 58.910 147.240 ;
        RECT 59.185 147.175 60.850 147.345 ;
        RECT 61.035 147.190 61.325 147.915 ;
        RECT 62.530 147.285 62.815 147.745 ;
        RECT 62.985 147.455 63.255 147.915 ;
        RECT 59.185 147.005 59.355 147.175 ;
        RECT 62.530 147.115 63.485 147.285 ;
        RECT 59.080 146.675 59.355 147.005 ;
        RECT 59.525 146.675 60.350 147.005 ;
        RECT 60.520 146.675 60.865 147.005 ;
        RECT 59.185 146.505 59.355 146.675 ;
        RECT 57.315 145.535 57.815 145.955 ;
        RECT 58.305 145.365 58.515 145.825 ;
        RECT 58.740 145.535 59.015 146.505 ;
        RECT 59.185 146.335 59.845 146.505 ;
        RECT 60.155 146.385 60.350 146.675 ;
        RECT 59.675 146.215 59.845 146.335 ;
        RECT 60.520 146.215 60.845 146.505 ;
        RECT 59.225 145.365 59.505 146.165 ;
        RECT 59.675 146.045 60.845 146.215 ;
        RECT 59.675 145.585 60.865 145.875 ;
        RECT 61.035 145.365 61.325 146.530 ;
        RECT 62.415 146.385 63.105 146.945 ;
        RECT 63.275 146.215 63.485 147.115 ;
        RECT 62.530 145.995 63.485 146.215 ;
        RECT 63.655 146.945 64.055 147.745 ;
        RECT 64.245 147.285 64.525 147.745 ;
        RECT 65.045 147.455 65.370 147.915 ;
        RECT 64.245 147.115 65.370 147.285 ;
        RECT 65.540 147.175 65.925 147.745 ;
        RECT 64.920 147.005 65.370 147.115 ;
        RECT 63.655 146.385 64.750 146.945 ;
        RECT 64.920 146.675 65.475 147.005 ;
        RECT 62.530 145.535 62.815 145.995 ;
        RECT 62.985 145.365 63.255 145.825 ;
        RECT 63.655 145.535 64.055 146.385 ;
        RECT 64.920 146.215 65.370 146.675 ;
        RECT 65.645 146.505 65.925 147.175 ;
        RECT 64.245 145.995 65.370 146.215 ;
        RECT 64.245 145.535 64.525 145.995 ;
        RECT 65.045 145.365 65.370 145.825 ;
        RECT 65.540 145.535 65.925 146.505 ;
        RECT 66.100 147.240 66.375 147.585 ;
        RECT 66.565 147.515 66.945 147.915 ;
        RECT 67.115 147.345 67.285 147.695 ;
        RECT 67.455 147.515 67.785 147.915 ;
        RECT 67.955 147.345 68.210 147.695 ;
        RECT 66.100 146.505 66.270 147.240 ;
        RECT 66.545 147.175 68.210 147.345 ;
        RECT 68.395 147.175 68.905 147.745 ;
        RECT 69.075 147.355 69.245 147.915 ;
        RECT 69.450 147.345 69.780 147.745 ;
        RECT 69.955 147.515 70.285 147.915 ;
        RECT 70.520 147.535 71.905 147.745 ;
        RECT 70.520 147.345 70.850 147.535 ;
        RECT 69.450 147.175 70.850 147.345 ;
        RECT 71.020 147.175 71.445 147.365 ;
        RECT 71.615 147.265 71.905 147.535 ;
        RECT 72.075 147.265 72.335 147.745 ;
        RECT 72.505 147.455 72.835 147.915 ;
        RECT 73.025 147.275 73.225 147.695 ;
        RECT 66.545 147.005 66.715 147.175 ;
        RECT 66.440 146.675 66.715 147.005 ;
        RECT 66.885 146.675 67.710 147.005 ;
        RECT 67.880 146.675 68.225 147.005 ;
        RECT 66.545 146.505 66.715 146.675 ;
        RECT 66.100 145.535 66.375 146.505 ;
        RECT 66.545 146.335 67.205 146.505 ;
        RECT 67.515 146.385 67.710 146.675 ;
        RECT 68.395 146.505 68.570 147.175 ;
        RECT 68.755 146.925 68.945 147.005 ;
        RECT 69.315 146.925 69.485 147.005 ;
        RECT 68.755 146.675 69.120 146.925 ;
        RECT 69.315 146.675 69.565 146.925 ;
        RECT 69.775 146.675 70.120 147.005 ;
        RECT 68.950 146.505 69.120 146.675 ;
        RECT 67.035 146.215 67.205 146.335 ;
        RECT 67.880 146.215 68.205 146.505 ;
        RECT 66.585 145.365 66.865 146.165 ;
        RECT 67.035 146.045 68.205 146.215 ;
        RECT 67.035 145.585 68.225 145.875 ;
        RECT 68.395 145.545 68.780 146.505 ;
        RECT 68.950 146.335 69.625 146.505 ;
        RECT 68.995 145.365 69.285 146.165 ;
        RECT 69.455 145.705 69.625 146.335 ;
        RECT 69.795 145.875 70.120 146.675 ;
        RECT 70.290 146.340 70.565 147.005 ;
        RECT 70.750 146.340 71.105 147.005 ;
        RECT 71.275 146.165 71.445 147.175 ;
        RECT 71.630 146.675 71.905 147.005 ;
        RECT 70.490 145.915 71.445 146.165 ;
        RECT 70.490 145.705 70.820 145.915 ;
        RECT 69.455 145.535 70.820 145.705 ;
        RECT 71.615 145.365 71.905 146.505 ;
        RECT 72.075 146.235 72.245 147.265 ;
        RECT 72.415 146.575 72.645 147.005 ;
        RECT 72.815 146.755 73.225 147.275 ;
        RECT 73.395 147.430 74.185 147.695 ;
        RECT 73.395 146.575 73.650 147.430 ;
        RECT 74.365 147.095 74.695 147.515 ;
        RECT 74.865 147.095 75.125 147.915 ;
        RECT 75.295 147.115 75.990 147.745 ;
        RECT 76.195 147.115 76.505 147.915 ;
        RECT 76.675 147.175 77.185 147.745 ;
        RECT 77.355 147.355 77.525 147.915 ;
        RECT 77.730 147.345 78.060 147.745 ;
        RECT 78.235 147.515 78.565 147.915 ;
        RECT 78.800 147.535 80.185 147.745 ;
        RECT 78.800 147.345 79.130 147.535 ;
        RECT 77.730 147.175 79.130 147.345 ;
        RECT 79.300 147.175 79.725 147.365 ;
        RECT 79.895 147.265 80.185 147.535 ;
        RECT 80.830 147.345 81.085 147.695 ;
        RECT 81.255 147.515 81.585 147.915 ;
        RECT 81.755 147.345 81.925 147.695 ;
        RECT 82.095 147.515 82.475 147.915 ;
        RECT 80.830 147.175 82.495 147.345 ;
        RECT 82.665 147.240 82.940 147.585 ;
        RECT 74.365 147.005 74.615 147.095 ;
        RECT 73.820 146.755 74.615 147.005 ;
        RECT 72.415 146.405 74.205 146.575 ;
        RECT 72.075 145.535 72.350 146.235 ;
        RECT 72.520 146.110 73.235 146.405 ;
        RECT 73.455 146.045 73.785 146.235 ;
        RECT 72.560 145.365 72.775 145.910 ;
        RECT 72.945 145.535 73.420 145.875 ;
        RECT 73.590 145.870 73.785 146.045 ;
        RECT 73.955 146.040 74.205 146.405 ;
        RECT 73.590 145.365 74.205 145.870 ;
        RECT 74.445 145.535 74.615 146.755 ;
        RECT 74.785 146.045 75.125 146.925 ;
        RECT 75.315 146.675 75.650 146.925 ;
        RECT 75.820 146.515 75.990 147.115 ;
        RECT 76.160 146.675 76.495 146.945 ;
        RECT 74.865 145.365 75.125 145.875 ;
        RECT 75.295 145.365 75.555 146.505 ;
        RECT 75.725 145.535 76.055 146.515 ;
        RECT 76.675 146.505 76.850 147.175 ;
        RECT 77.035 146.925 77.225 147.005 ;
        RECT 77.595 146.925 77.765 147.005 ;
        RECT 77.035 146.675 77.400 146.925 ;
        RECT 77.595 146.675 77.845 146.925 ;
        RECT 78.055 146.675 78.400 147.005 ;
        RECT 77.230 146.505 77.400 146.675 ;
        RECT 76.225 145.365 76.505 146.505 ;
        RECT 76.675 145.545 77.060 146.505 ;
        RECT 77.230 146.335 77.905 146.505 ;
        RECT 77.275 145.365 77.565 146.165 ;
        RECT 77.735 145.705 77.905 146.335 ;
        RECT 78.075 145.875 78.400 146.675 ;
        RECT 78.570 146.340 78.845 147.005 ;
        RECT 79.030 146.340 79.385 147.005 ;
        RECT 79.555 146.165 79.725 147.175 ;
        RECT 82.325 147.005 82.495 147.175 ;
        RECT 79.910 146.675 80.185 147.005 ;
        RECT 80.815 146.675 81.160 147.005 ;
        RECT 81.330 146.675 82.155 147.005 ;
        RECT 82.325 146.675 82.600 147.005 ;
        RECT 78.770 145.915 79.725 146.165 ;
        RECT 78.770 145.705 79.100 145.915 ;
        RECT 77.735 145.535 79.100 145.705 ;
        RECT 79.895 145.365 80.185 146.505 ;
        RECT 80.835 146.215 81.160 146.505 ;
        RECT 81.330 146.385 81.525 146.675 ;
        RECT 82.325 146.505 82.495 146.675 ;
        RECT 82.770 146.505 82.940 147.240 ;
        RECT 83.120 147.385 83.410 147.735 ;
        RECT 83.605 147.555 83.935 147.915 ;
        RECT 84.105 147.385 84.335 147.690 ;
        RECT 83.120 147.215 84.335 147.385 ;
        RECT 84.525 147.235 84.695 147.610 ;
        RECT 84.525 147.065 84.725 147.235 ;
        RECT 84.965 147.105 85.235 147.915 ;
        RECT 85.405 147.105 85.735 147.745 ;
        RECT 85.905 147.105 86.145 147.915 ;
        RECT 86.795 147.190 87.085 147.915 ;
        RECT 87.260 147.150 87.715 147.915 ;
        RECT 87.990 147.535 89.290 147.745 ;
        RECT 89.545 147.555 89.875 147.915 ;
        RECT 89.120 147.385 89.290 147.535 ;
        RECT 90.045 147.415 90.305 147.745 ;
        RECT 90.075 147.405 90.305 147.415 ;
        RECT 84.525 147.045 84.695 147.065 ;
        RECT 83.180 146.895 83.440 147.005 ;
        RECT 83.175 146.725 83.440 146.895 ;
        RECT 83.180 146.675 83.440 146.725 ;
        RECT 83.620 146.675 84.005 147.005 ;
        RECT 84.175 146.875 84.695 147.045 ;
        RECT 81.835 146.335 82.495 146.505 ;
        RECT 81.835 146.215 82.005 146.335 ;
        RECT 80.835 146.045 82.005 146.215 ;
        RECT 80.815 145.585 82.005 145.875 ;
        RECT 82.175 145.365 82.455 146.165 ;
        RECT 82.665 145.535 82.940 146.505 ;
        RECT 83.120 145.365 83.440 146.505 ;
        RECT 83.620 145.625 83.815 146.675 ;
        RECT 84.175 146.495 84.345 146.875 ;
        RECT 83.995 146.215 84.345 146.495 ;
        RECT 84.535 146.345 84.780 146.705 ;
        RECT 84.955 146.675 85.305 146.925 ;
        RECT 85.475 146.505 85.645 147.105 ;
        RECT 88.190 146.925 88.410 147.325 ;
        RECT 85.815 146.675 86.165 146.925 ;
        RECT 87.255 146.725 87.745 146.925 ;
        RECT 87.935 146.715 88.410 146.925 ;
        RECT 88.655 146.925 88.865 147.325 ;
        RECT 89.120 147.260 89.875 147.385 ;
        RECT 89.120 147.215 89.965 147.260 ;
        RECT 89.695 147.095 89.965 147.215 ;
        RECT 88.655 146.715 88.985 146.925 ;
        RECT 89.155 146.655 89.565 146.960 ;
        RECT 83.995 145.535 84.325 146.215 ;
        RECT 84.525 145.365 84.780 146.165 ;
        RECT 84.965 145.365 85.295 146.505 ;
        RECT 85.475 146.335 86.155 146.505 ;
        RECT 85.825 145.550 86.155 146.335 ;
        RECT 86.795 145.365 87.085 146.530 ;
        RECT 87.260 146.485 88.435 146.545 ;
        RECT 89.795 146.520 89.965 147.095 ;
        RECT 89.765 146.485 89.965 146.520 ;
        RECT 87.260 146.375 89.965 146.485 ;
        RECT 87.260 145.755 87.515 146.375 ;
        RECT 88.105 146.315 89.905 146.375 ;
        RECT 88.105 146.285 88.435 146.315 ;
        RECT 90.135 146.215 90.305 147.405 ;
        RECT 90.475 147.370 95.820 147.915 ;
        RECT 95.995 147.370 101.340 147.915 ;
        RECT 101.515 147.370 106.860 147.915 ;
        RECT 92.060 146.540 92.400 147.370 ;
        RECT 87.765 146.115 87.950 146.205 ;
        RECT 88.540 146.115 89.375 146.125 ;
        RECT 87.765 145.915 89.375 146.115 ;
        RECT 87.765 145.875 87.995 145.915 ;
        RECT 87.260 145.535 87.595 145.755 ;
        RECT 88.600 145.365 88.955 145.745 ;
        RECT 89.125 145.535 89.375 145.915 ;
        RECT 89.625 145.365 89.875 146.145 ;
        RECT 90.045 145.535 90.305 146.215 ;
        RECT 93.880 145.800 94.230 147.050 ;
        RECT 97.580 146.540 97.920 147.370 ;
        RECT 99.400 145.800 99.750 147.050 ;
        RECT 103.100 146.540 103.440 147.370 ;
        RECT 107.955 147.165 109.165 147.915 ;
        RECT 104.920 145.800 105.270 147.050 ;
        RECT 107.955 146.455 108.475 146.995 ;
        RECT 108.645 146.625 109.165 147.165 ;
        RECT 90.475 145.365 95.820 145.800 ;
        RECT 95.995 145.365 101.340 145.800 ;
        RECT 101.515 145.365 106.860 145.800 ;
        RECT 107.955 145.365 109.165 146.455 ;
        RECT 35.190 145.195 109.250 145.365 ;
        RECT 35.275 144.105 36.485 145.195 ;
        RECT 36.655 144.760 42.000 145.195 ;
        RECT 42.175 144.760 47.520 145.195 ;
        RECT 35.275 143.395 35.795 143.935 ;
        RECT 35.965 143.565 36.485 144.105 ;
        RECT 35.275 142.645 36.485 143.395 ;
        RECT 38.240 143.190 38.580 144.020 ;
        RECT 40.060 143.510 40.410 144.760 ;
        RECT 43.760 143.190 44.100 144.020 ;
        RECT 45.580 143.510 45.930 144.760 ;
        RECT 48.155 144.030 48.445 145.195 ;
        RECT 48.615 144.760 53.960 145.195 ;
        RECT 36.655 142.645 42.000 143.190 ;
        RECT 42.175 142.645 47.520 143.190 ;
        RECT 48.155 142.645 48.445 143.370 ;
        RECT 50.200 143.190 50.540 144.020 ;
        RECT 52.020 143.510 52.370 144.760 ;
        RECT 55.145 144.450 55.415 145.195 ;
        RECT 56.045 145.190 62.320 145.195 ;
        RECT 55.585 144.280 55.875 145.020 ;
        RECT 56.045 144.465 56.300 145.190 ;
        RECT 56.485 144.295 56.745 145.020 ;
        RECT 56.915 144.465 57.160 145.190 ;
        RECT 57.345 144.295 57.605 145.020 ;
        RECT 57.775 144.465 58.020 145.190 ;
        RECT 58.205 144.295 58.465 145.020 ;
        RECT 58.635 144.465 58.880 145.190 ;
        RECT 59.050 144.295 59.310 145.020 ;
        RECT 59.480 144.465 59.740 145.190 ;
        RECT 59.910 144.295 60.170 145.020 ;
        RECT 60.340 144.465 60.600 145.190 ;
        RECT 60.770 144.295 61.030 145.020 ;
        RECT 61.200 144.465 61.460 145.190 ;
        RECT 61.630 144.295 61.890 145.020 ;
        RECT 62.060 144.395 62.320 145.190 ;
        RECT 56.485 144.280 61.890 144.295 ;
        RECT 55.145 144.055 61.890 144.280 ;
        RECT 55.145 143.465 56.310 144.055 ;
        RECT 62.490 143.885 62.740 145.020 ;
        RECT 62.920 144.385 63.180 145.195 ;
        RECT 63.355 143.885 63.600 145.025 ;
        RECT 63.780 144.385 64.075 145.195 ;
        RECT 64.725 144.385 65.020 145.195 ;
        RECT 65.200 143.885 65.445 145.025 ;
        RECT 65.620 144.385 65.880 145.195 ;
        RECT 66.480 145.190 72.755 145.195 ;
        RECT 66.060 143.885 66.310 145.020 ;
        RECT 66.480 144.395 66.740 145.190 ;
        RECT 66.910 144.295 67.170 145.020 ;
        RECT 67.340 144.465 67.600 145.190 ;
        RECT 67.770 144.295 68.030 145.020 ;
        RECT 68.200 144.465 68.460 145.190 ;
        RECT 68.630 144.295 68.890 145.020 ;
        RECT 69.060 144.465 69.320 145.190 ;
        RECT 69.490 144.295 69.750 145.020 ;
        RECT 69.920 144.465 70.165 145.190 ;
        RECT 70.335 144.295 70.595 145.020 ;
        RECT 70.780 144.465 71.025 145.190 ;
        RECT 71.195 144.295 71.455 145.020 ;
        RECT 71.640 144.465 71.885 145.190 ;
        RECT 72.055 144.295 72.315 145.020 ;
        RECT 72.500 144.465 72.755 145.190 ;
        RECT 66.910 144.280 72.315 144.295 ;
        RECT 72.925 144.280 73.215 145.020 ;
        RECT 73.385 144.450 73.655 145.195 ;
        RECT 66.910 144.055 73.655 144.280 ;
        RECT 56.480 143.635 63.600 143.885 ;
        RECT 55.145 143.295 61.890 143.465 ;
        RECT 48.615 142.645 53.960 143.190 ;
        RECT 55.145 142.645 55.445 143.125 ;
        RECT 55.615 142.840 55.875 143.295 ;
        RECT 56.045 142.645 56.305 143.125 ;
        RECT 56.485 142.840 56.745 143.295 ;
        RECT 56.915 142.645 57.165 143.125 ;
        RECT 57.345 142.840 57.605 143.295 ;
        RECT 57.775 142.645 58.025 143.125 ;
        RECT 58.205 142.840 58.465 143.295 ;
        RECT 58.635 142.645 58.880 143.125 ;
        RECT 59.050 142.840 59.325 143.295 ;
        RECT 59.495 142.645 59.740 143.125 ;
        RECT 59.910 142.840 60.170 143.295 ;
        RECT 60.340 142.645 60.600 143.125 ;
        RECT 60.770 142.840 61.030 143.295 ;
        RECT 61.200 142.645 61.460 143.125 ;
        RECT 61.630 142.840 61.890 143.295 ;
        RECT 62.060 142.645 62.320 143.205 ;
        RECT 62.490 142.825 62.740 143.635 ;
        RECT 62.920 142.645 63.180 143.170 ;
        RECT 63.350 142.825 63.600 143.635 ;
        RECT 63.770 143.325 64.085 143.885 ;
        RECT 64.715 143.325 65.030 143.885 ;
        RECT 65.200 143.635 72.320 143.885 ;
        RECT 63.780 142.645 64.085 143.155 ;
        RECT 64.715 142.645 65.020 143.155 ;
        RECT 65.200 142.825 65.450 143.635 ;
        RECT 65.620 142.645 65.880 143.170 ;
        RECT 66.060 142.825 66.310 143.635 ;
        RECT 72.490 143.495 73.655 144.055 ;
        RECT 73.915 144.030 74.205 145.195 ;
        RECT 74.400 144.225 74.700 144.420 ;
        RECT 74.870 144.395 75.125 145.195 ;
        RECT 75.325 144.565 75.655 145.025 ;
        RECT 75.825 144.735 76.400 145.195 ;
        RECT 76.570 144.565 76.925 145.025 ;
        RECT 75.325 144.395 76.925 144.565 ;
        RECT 74.400 144.055 75.650 144.225 ;
        RECT 72.490 143.465 73.685 143.495 ;
        RECT 66.910 143.325 73.685 143.465 ;
        RECT 74.400 143.400 74.570 144.055 ;
        RECT 74.745 143.555 75.090 143.885 ;
        RECT 75.320 143.635 75.650 144.055 ;
        RECT 75.820 143.495 76.100 144.395 ;
        RECT 76.280 143.835 76.470 144.215 ;
        RECT 76.650 144.055 76.925 144.395 ;
        RECT 77.095 144.055 77.425 145.195 ;
        RECT 77.595 144.105 81.105 145.195 ;
        RECT 76.280 143.635 77.425 143.835 ;
        RECT 75.815 143.465 76.100 143.495 ;
        RECT 66.910 143.295 73.655 143.325 ;
        RECT 66.480 142.645 66.740 143.205 ;
        RECT 66.910 142.840 67.170 143.295 ;
        RECT 67.340 142.645 67.600 143.125 ;
        RECT 67.770 142.840 68.030 143.295 ;
        RECT 68.200 142.645 68.460 143.125 ;
        RECT 68.630 142.840 68.890 143.295 ;
        RECT 69.060 142.645 69.305 143.125 ;
        RECT 69.475 142.840 69.750 143.295 ;
        RECT 69.920 142.645 70.165 143.125 ;
        RECT 70.335 142.840 70.595 143.295 ;
        RECT 70.775 142.645 71.025 143.125 ;
        RECT 71.195 142.840 71.455 143.295 ;
        RECT 71.635 142.645 71.885 143.125 ;
        RECT 72.055 142.840 72.315 143.295 ;
        RECT 72.495 142.645 72.755 143.125 ;
        RECT 72.925 142.840 73.185 143.295 ;
        RECT 73.355 142.645 73.655 143.125 ;
        RECT 73.915 142.645 74.205 143.370 ;
        RECT 74.400 143.070 74.635 143.400 ;
        RECT 74.805 142.645 75.135 143.385 ;
        RECT 75.370 143.025 75.645 143.465 ;
        RECT 75.815 143.195 76.145 143.465 ;
        RECT 76.315 143.255 77.425 143.465 ;
        RECT 76.315 143.025 76.565 143.255 ;
        RECT 75.370 142.815 76.565 143.025 ;
        RECT 76.735 142.645 76.905 143.085 ;
        RECT 77.075 142.815 77.425 143.255 ;
        RECT 77.595 143.415 79.245 143.935 ;
        RECT 79.415 143.585 81.105 144.105 ;
        RECT 82.235 144.055 82.465 145.195 ;
        RECT 82.635 144.045 82.965 145.025 ;
        RECT 83.135 144.055 83.345 145.195 ;
        RECT 83.575 144.760 88.920 145.195 ;
        RECT 89.095 144.760 94.440 145.195 ;
        RECT 82.215 143.635 82.545 143.885 ;
        RECT 77.595 142.645 81.105 143.415 ;
        RECT 82.235 142.645 82.465 143.465 ;
        RECT 82.715 143.445 82.965 144.045 ;
        RECT 82.635 142.815 82.965 143.445 ;
        RECT 83.135 142.645 83.345 143.465 ;
        RECT 85.160 143.190 85.500 144.020 ;
        RECT 86.980 143.510 87.330 144.760 ;
        RECT 90.680 143.190 91.020 144.020 ;
        RECT 92.500 143.510 92.850 144.760 ;
        RECT 94.615 144.105 95.825 145.195 ;
        RECT 94.615 143.395 95.135 143.935 ;
        RECT 95.305 143.565 95.825 144.105 ;
        RECT 96.035 144.055 96.265 145.195 ;
        RECT 96.435 144.045 96.765 145.025 ;
        RECT 96.935 144.055 97.145 145.195 ;
        RECT 97.375 144.105 99.045 145.195 ;
        RECT 96.015 143.635 96.345 143.885 ;
        RECT 83.575 142.645 88.920 143.190 ;
        RECT 89.095 142.645 94.440 143.190 ;
        RECT 94.615 142.645 95.825 143.395 ;
        RECT 96.035 142.645 96.265 143.465 ;
        RECT 96.515 143.445 96.765 144.045 ;
        RECT 96.435 142.815 96.765 143.445 ;
        RECT 96.935 142.645 97.145 143.465 ;
        RECT 97.375 143.415 98.125 143.935 ;
        RECT 98.295 143.585 99.045 144.105 ;
        RECT 99.675 144.030 99.965 145.195 ;
        RECT 100.135 144.760 105.480 145.195 ;
        RECT 97.375 142.645 99.045 143.415 ;
        RECT 99.675 142.645 99.965 143.370 ;
        RECT 101.720 143.190 102.060 144.020 ;
        RECT 103.540 143.510 103.890 144.760 ;
        RECT 105.655 144.105 107.325 145.195 ;
        RECT 105.655 143.415 106.405 143.935 ;
        RECT 106.575 143.585 107.325 144.105 ;
        RECT 107.955 144.105 109.165 145.195 ;
        RECT 107.955 143.565 108.475 144.105 ;
        RECT 100.135 142.645 105.480 143.190 ;
        RECT 105.655 142.645 107.325 143.415 ;
        RECT 108.645 143.395 109.165 143.935 ;
        RECT 107.955 142.645 109.165 143.395 ;
        RECT 35.190 142.475 109.250 142.645 ;
        RECT 35.275 141.725 36.485 142.475 ;
        RECT 36.655 141.930 42.000 142.475 ;
        RECT 35.275 141.185 35.795 141.725 ;
        RECT 35.965 141.015 36.485 141.555 ;
        RECT 38.240 141.100 38.580 141.930 ;
        RECT 42.640 141.925 42.895 142.215 ;
        RECT 43.065 142.095 43.395 142.475 ;
        RECT 42.640 141.755 43.390 141.925 ;
        RECT 35.275 139.925 36.485 141.015 ;
        RECT 40.060 140.360 40.410 141.610 ;
        RECT 42.640 140.935 42.990 141.585 ;
        RECT 43.160 140.765 43.390 141.755 ;
        RECT 42.640 140.595 43.390 140.765 ;
        RECT 36.655 139.925 42.000 140.360 ;
        RECT 42.640 140.095 42.895 140.595 ;
        RECT 43.065 139.925 43.395 140.425 ;
        RECT 43.565 140.095 43.735 142.215 ;
        RECT 44.095 142.115 44.425 142.475 ;
        RECT 44.595 142.085 45.090 142.255 ;
        RECT 45.295 142.085 46.150 142.255 ;
        RECT 43.965 140.895 44.425 141.945 ;
        RECT 43.905 140.110 44.230 140.895 ;
        RECT 44.595 140.725 44.765 142.085 ;
        RECT 44.935 141.175 45.285 141.795 ;
        RECT 45.455 141.575 45.810 141.795 ;
        RECT 45.455 140.985 45.625 141.575 ;
        RECT 45.980 141.375 46.150 142.085 ;
        RECT 47.025 142.015 47.355 142.475 ;
        RECT 47.565 142.115 47.915 142.285 ;
        RECT 46.355 141.545 47.145 141.795 ;
        RECT 47.565 141.725 47.825 142.115 ;
        RECT 48.135 142.025 49.085 142.305 ;
        RECT 49.255 142.035 49.445 142.475 ;
        RECT 49.615 142.095 50.685 142.265 ;
        RECT 47.315 141.375 47.485 141.555 ;
        RECT 44.595 140.555 44.990 140.725 ;
        RECT 45.160 140.595 45.625 140.985 ;
        RECT 45.795 141.205 47.485 141.375 ;
        RECT 44.820 140.425 44.990 140.555 ;
        RECT 45.795 140.425 45.965 141.205 ;
        RECT 47.655 141.035 47.825 141.725 ;
        RECT 46.325 140.865 47.825 141.035 ;
        RECT 48.015 141.065 48.225 141.855 ;
        RECT 48.395 141.235 48.745 141.855 ;
        RECT 48.915 141.245 49.085 142.025 ;
        RECT 49.615 141.865 49.785 142.095 ;
        RECT 49.255 141.695 49.785 141.865 ;
        RECT 49.255 141.415 49.475 141.695 ;
        RECT 49.955 141.525 50.195 141.925 ;
        RECT 48.915 141.075 49.320 141.245 ;
        RECT 49.655 141.155 50.195 141.525 ;
        RECT 50.365 141.740 50.685 142.095 ;
        RECT 50.930 142.015 51.235 142.475 ;
        RECT 51.405 141.765 51.660 142.295 ;
        RECT 50.365 141.565 50.690 141.740 ;
        RECT 50.365 141.265 51.280 141.565 ;
        RECT 50.540 141.235 51.280 141.265 ;
        RECT 48.015 140.905 48.690 141.065 ;
        RECT 49.150 140.985 49.320 141.075 ;
        RECT 48.015 140.895 48.980 140.905 ;
        RECT 47.655 140.725 47.825 140.865 ;
        RECT 44.400 139.925 44.650 140.385 ;
        RECT 44.820 140.095 45.070 140.425 ;
        RECT 45.285 140.095 45.965 140.425 ;
        RECT 46.135 140.525 47.210 140.695 ;
        RECT 47.655 140.555 48.215 140.725 ;
        RECT 48.520 140.605 48.980 140.895 ;
        RECT 49.150 140.815 50.370 140.985 ;
        RECT 46.135 140.185 46.305 140.525 ;
        RECT 46.540 139.925 46.870 140.355 ;
        RECT 47.040 140.185 47.210 140.525 ;
        RECT 47.505 139.925 47.875 140.385 ;
        RECT 48.045 140.095 48.215 140.555 ;
        RECT 49.150 140.435 49.320 140.815 ;
        RECT 50.540 140.645 50.710 141.235 ;
        RECT 51.450 141.115 51.660 141.765 ;
        RECT 51.840 141.925 52.095 142.215 ;
        RECT 52.265 142.095 52.595 142.475 ;
        RECT 51.840 141.755 52.590 141.925 ;
        RECT 48.450 140.095 49.320 140.435 ;
        RECT 49.910 140.475 50.710 140.645 ;
        RECT 49.490 139.925 49.740 140.385 ;
        RECT 49.910 140.185 50.080 140.475 ;
        RECT 50.260 139.925 50.590 140.305 ;
        RECT 50.930 139.925 51.235 141.065 ;
        RECT 51.405 140.235 51.660 141.115 ;
        RECT 51.840 140.935 52.190 141.585 ;
        RECT 52.360 140.765 52.590 141.755 ;
        RECT 51.840 140.595 52.590 140.765 ;
        RECT 51.840 140.095 52.095 140.595 ;
        RECT 52.265 139.925 52.595 140.425 ;
        RECT 52.765 140.095 52.935 142.215 ;
        RECT 53.295 142.115 53.625 142.475 ;
        RECT 53.795 142.085 54.290 142.255 ;
        RECT 54.495 142.085 55.350 142.255 ;
        RECT 53.165 140.895 53.625 141.945 ;
        RECT 53.105 140.110 53.430 140.895 ;
        RECT 53.795 140.725 53.965 142.085 ;
        RECT 54.135 141.175 54.485 141.795 ;
        RECT 54.655 141.575 55.010 141.795 ;
        RECT 54.655 140.985 54.825 141.575 ;
        RECT 55.180 141.375 55.350 142.085 ;
        RECT 56.225 142.015 56.555 142.475 ;
        RECT 56.765 142.115 57.115 142.285 ;
        RECT 55.555 141.545 56.345 141.795 ;
        RECT 56.765 141.725 57.025 142.115 ;
        RECT 57.335 142.025 58.285 142.305 ;
        RECT 58.455 142.035 58.645 142.475 ;
        RECT 58.815 142.095 59.885 142.265 ;
        RECT 56.515 141.375 56.685 141.555 ;
        RECT 53.795 140.555 54.190 140.725 ;
        RECT 54.360 140.595 54.825 140.985 ;
        RECT 54.995 141.205 56.685 141.375 ;
        RECT 54.020 140.425 54.190 140.555 ;
        RECT 54.995 140.425 55.165 141.205 ;
        RECT 56.855 141.035 57.025 141.725 ;
        RECT 55.525 140.865 57.025 141.035 ;
        RECT 57.215 141.065 57.425 141.855 ;
        RECT 57.595 141.235 57.945 141.855 ;
        RECT 58.115 141.245 58.285 142.025 ;
        RECT 58.815 141.865 58.985 142.095 ;
        RECT 58.455 141.695 58.985 141.865 ;
        RECT 58.455 141.415 58.675 141.695 ;
        RECT 59.155 141.525 59.395 141.925 ;
        RECT 58.115 141.075 58.520 141.245 ;
        RECT 58.855 141.155 59.395 141.525 ;
        RECT 59.565 141.740 59.885 142.095 ;
        RECT 60.130 142.015 60.435 142.475 ;
        RECT 60.605 141.765 60.860 142.295 ;
        RECT 59.565 141.565 59.890 141.740 ;
        RECT 59.565 141.265 60.480 141.565 ;
        RECT 59.740 141.235 60.480 141.265 ;
        RECT 57.215 140.905 57.890 141.065 ;
        RECT 58.350 140.985 58.520 141.075 ;
        RECT 57.215 140.895 58.180 140.905 ;
        RECT 56.855 140.725 57.025 140.865 ;
        RECT 53.600 139.925 53.850 140.385 ;
        RECT 54.020 140.095 54.270 140.425 ;
        RECT 54.485 140.095 55.165 140.425 ;
        RECT 55.335 140.525 56.410 140.695 ;
        RECT 56.855 140.555 57.415 140.725 ;
        RECT 57.720 140.605 58.180 140.895 ;
        RECT 58.350 140.815 59.570 140.985 ;
        RECT 55.335 140.185 55.505 140.525 ;
        RECT 55.740 139.925 56.070 140.355 ;
        RECT 56.240 140.185 56.410 140.525 ;
        RECT 56.705 139.925 57.075 140.385 ;
        RECT 57.245 140.095 57.415 140.555 ;
        RECT 58.350 140.435 58.520 140.815 ;
        RECT 59.740 140.645 59.910 141.235 ;
        RECT 60.650 141.115 60.860 141.765 ;
        RECT 61.035 141.750 61.325 142.475 ;
        RECT 61.495 141.750 61.755 142.305 ;
        RECT 61.925 142.030 62.355 142.475 ;
        RECT 62.590 141.905 62.760 142.305 ;
        RECT 62.930 142.075 63.650 142.475 ;
        RECT 57.650 140.095 58.520 140.435 ;
        RECT 59.110 140.475 59.910 140.645 ;
        RECT 58.690 139.925 58.940 140.385 ;
        RECT 59.110 140.185 59.280 140.475 ;
        RECT 59.460 139.925 59.790 140.305 ;
        RECT 60.130 139.925 60.435 141.065 ;
        RECT 60.605 140.235 60.860 141.115 ;
        RECT 61.035 139.925 61.325 141.090 ;
        RECT 61.495 141.035 61.670 141.750 ;
        RECT 62.590 141.735 63.470 141.905 ;
        RECT 63.820 141.860 63.990 142.305 ;
        RECT 64.565 141.965 64.965 142.475 ;
        RECT 61.840 141.235 62.095 141.565 ;
        RECT 61.495 140.095 61.755 141.035 ;
        RECT 61.925 140.755 62.095 141.235 ;
        RECT 62.320 140.945 62.650 141.565 ;
        RECT 62.820 141.185 63.110 141.565 ;
        RECT 63.300 141.015 63.470 141.735 ;
        RECT 62.950 140.845 63.470 141.015 ;
        RECT 63.640 141.690 63.990 141.860 ;
        RECT 61.925 140.585 62.685 140.755 ;
        RECT 62.950 140.655 63.120 140.845 ;
        RECT 63.640 140.665 63.810 141.690 ;
        RECT 64.230 141.205 64.490 141.795 ;
        RECT 64.010 140.905 64.490 141.205 ;
        RECT 64.690 140.905 64.950 141.795 ;
        RECT 66.095 141.675 66.790 142.305 ;
        RECT 66.995 141.675 67.305 142.475 ;
        RECT 67.475 141.705 70.985 142.475 ;
        RECT 71.180 141.825 71.490 142.295 ;
        RECT 71.660 141.995 72.395 142.475 ;
        RECT 72.565 141.905 72.735 142.255 ;
        RECT 72.905 142.075 73.285 142.475 ;
        RECT 66.115 141.235 66.450 141.485 ;
        RECT 66.620 141.075 66.790 141.675 ;
        RECT 66.960 141.235 67.295 141.505 ;
        RECT 67.475 141.185 69.125 141.705 ;
        RECT 71.180 141.655 71.915 141.825 ;
        RECT 72.565 141.735 73.305 141.905 ;
        RECT 73.475 141.800 73.745 142.145 ;
        RECT 71.665 141.565 71.915 141.655 ;
        RECT 73.135 141.565 73.305 141.735 ;
        RECT 62.515 140.360 62.685 140.585 ;
        RECT 63.400 140.495 63.810 140.665 ;
        RECT 63.985 140.555 64.925 140.725 ;
        RECT 63.400 140.360 63.655 140.495 ;
        RECT 61.925 139.925 62.255 140.325 ;
        RECT 62.515 140.190 63.655 140.360 ;
        RECT 63.985 140.305 64.155 140.555 ;
        RECT 63.400 140.095 63.655 140.190 ;
        RECT 63.825 140.135 64.155 140.305 ;
        RECT 64.325 139.925 64.575 140.385 ;
        RECT 64.745 140.095 64.925 140.555 ;
        RECT 66.095 139.925 66.355 141.065 ;
        RECT 66.525 140.095 66.855 141.075 ;
        RECT 67.025 139.925 67.305 141.065 ;
        RECT 69.295 141.015 70.985 141.535 ;
        RECT 71.160 141.235 71.495 141.485 ;
        RECT 71.665 141.235 72.405 141.565 ;
        RECT 73.135 141.235 73.365 141.565 ;
        RECT 67.475 139.925 70.985 141.015 ;
        RECT 71.160 139.925 71.415 141.065 ;
        RECT 71.665 140.675 71.835 141.235 ;
        RECT 73.135 141.065 73.305 141.235 ;
        RECT 73.575 141.065 73.745 141.800 ;
        RECT 73.925 141.665 74.195 142.475 ;
        RECT 74.365 141.665 74.695 142.305 ;
        RECT 74.865 141.665 75.105 142.475 ;
        RECT 73.915 141.235 74.265 141.485 ;
        RECT 74.435 141.065 74.605 141.665 ;
        RECT 75.795 141.655 76.025 142.475 ;
        RECT 76.195 141.675 76.525 142.305 ;
        RECT 74.775 141.235 75.125 141.485 ;
        RECT 75.775 141.235 76.105 141.485 ;
        RECT 76.275 141.075 76.525 141.675 ;
        RECT 76.695 141.655 76.905 142.475 ;
        RECT 77.135 141.725 78.345 142.475 ;
        RECT 77.135 141.185 77.655 141.725 ;
        RECT 78.515 141.655 78.775 142.475 ;
        RECT 78.945 141.655 79.275 142.075 ;
        RECT 79.455 141.905 79.715 142.305 ;
        RECT 79.885 142.075 80.215 142.475 ;
        RECT 80.385 141.905 80.555 142.255 ;
        RECT 80.725 142.075 81.100 142.475 ;
        RECT 79.455 141.735 81.120 141.905 ;
        RECT 81.290 141.800 81.565 142.145 ;
        RECT 79.025 141.565 79.275 141.655 ;
        RECT 80.950 141.565 81.120 141.735 ;
        RECT 72.060 140.895 73.305 141.065 ;
        RECT 72.060 140.645 72.480 140.895 ;
        RECT 71.610 140.145 72.805 140.475 ;
        RECT 72.985 139.925 73.265 140.725 ;
        RECT 73.475 140.095 73.745 141.065 ;
        RECT 73.925 139.925 74.255 141.065 ;
        RECT 74.435 140.895 75.115 141.065 ;
        RECT 74.785 140.110 75.115 140.895 ;
        RECT 75.795 139.925 76.025 141.065 ;
        RECT 76.195 140.095 76.525 141.075 ;
        RECT 76.695 139.925 76.905 141.065 ;
        RECT 77.825 141.015 78.345 141.555 ;
        RECT 78.520 141.235 78.855 141.485 ;
        RECT 79.025 141.235 79.740 141.565 ;
        RECT 79.955 141.235 80.780 141.565 ;
        RECT 80.950 141.235 81.225 141.565 ;
        RECT 77.135 139.925 78.345 141.015 ;
        RECT 78.515 139.925 78.775 141.065 ;
        RECT 79.025 140.675 79.195 141.235 ;
        RECT 79.455 140.775 79.785 141.065 ;
        RECT 79.955 140.945 80.200 141.235 ;
        RECT 80.950 141.065 81.120 141.235 ;
        RECT 81.395 141.065 81.565 141.800 ;
        RECT 82.665 141.755 82.995 142.475 ;
        RECT 83.540 142.075 85.155 142.245 ;
        RECT 85.325 142.075 85.655 142.475 ;
        RECT 84.985 141.905 85.155 142.075 ;
        RECT 85.825 142.000 86.160 142.260 ;
        RECT 82.720 141.235 83.070 141.565 ;
        RECT 83.380 141.235 83.800 141.900 ;
        RECT 83.970 141.455 84.260 141.895 ;
        RECT 84.450 141.795 84.720 141.895 ;
        RECT 84.450 141.625 84.725 141.795 ;
        RECT 84.985 141.735 85.545 141.905 ;
        RECT 83.970 141.285 84.265 141.455 ;
        RECT 83.970 141.235 84.260 141.285 ;
        RECT 84.450 141.235 84.720 141.625 ;
        RECT 85.375 141.565 85.545 141.735 ;
        RECT 84.930 141.455 85.180 141.565 ;
        RECT 84.930 141.285 85.185 141.455 ;
        RECT 84.930 141.235 85.180 141.285 ;
        RECT 85.375 141.235 85.680 141.565 ;
        RECT 82.720 141.115 82.925 141.235 ;
        RECT 80.460 140.895 81.120 141.065 ;
        RECT 80.460 140.775 80.630 140.895 ;
        RECT 79.455 140.605 80.630 140.775 ;
        RECT 79.015 140.105 80.630 140.435 ;
        RECT 80.800 139.925 81.080 140.725 ;
        RECT 81.290 140.095 81.565 141.065 ;
        RECT 82.715 140.945 82.925 141.115 ;
        RECT 85.375 141.065 85.545 141.235 ;
        RECT 83.175 140.895 85.545 141.065 ;
        RECT 82.745 140.265 82.915 140.765 ;
        RECT 83.175 140.435 83.345 140.895 ;
        RECT 83.575 140.515 85.000 140.685 ;
        RECT 83.575 140.265 83.905 140.515 ;
        RECT 82.745 140.095 83.905 140.265 ;
        RECT 84.130 139.925 84.460 140.345 ;
        RECT 84.715 140.095 85.000 140.515 ;
        RECT 85.245 139.925 85.575 140.725 ;
        RECT 85.905 140.645 86.160 142.000 ;
        RECT 86.795 141.750 87.085 142.475 ;
        RECT 87.260 141.925 87.515 142.215 ;
        RECT 87.685 142.095 88.015 142.475 ;
        RECT 87.260 141.755 88.010 141.925 ;
        RECT 85.825 140.135 86.160 140.645 ;
        RECT 86.795 139.925 87.085 141.090 ;
        RECT 87.260 140.935 87.610 141.585 ;
        RECT 87.780 140.765 88.010 141.755 ;
        RECT 87.260 140.595 88.010 140.765 ;
        RECT 87.260 140.095 87.515 140.595 ;
        RECT 87.685 139.925 88.015 140.425 ;
        RECT 88.185 140.095 88.355 142.215 ;
        RECT 88.715 142.115 89.045 142.475 ;
        RECT 89.215 142.085 89.710 142.255 ;
        RECT 89.915 142.085 90.770 142.255 ;
        RECT 88.585 140.895 89.045 141.945 ;
        RECT 88.525 140.110 88.850 140.895 ;
        RECT 89.215 140.725 89.385 142.085 ;
        RECT 89.555 141.175 89.905 141.795 ;
        RECT 90.075 141.575 90.430 141.795 ;
        RECT 90.075 140.985 90.245 141.575 ;
        RECT 90.600 141.375 90.770 142.085 ;
        RECT 91.645 142.015 91.975 142.475 ;
        RECT 92.185 142.115 92.535 142.285 ;
        RECT 90.975 141.545 91.765 141.795 ;
        RECT 92.185 141.725 92.445 142.115 ;
        RECT 92.755 142.025 93.705 142.305 ;
        RECT 93.875 142.035 94.065 142.475 ;
        RECT 94.235 142.095 95.305 142.265 ;
        RECT 91.935 141.375 92.105 141.555 ;
        RECT 89.215 140.555 89.610 140.725 ;
        RECT 89.780 140.595 90.245 140.985 ;
        RECT 90.415 141.205 92.105 141.375 ;
        RECT 89.440 140.425 89.610 140.555 ;
        RECT 90.415 140.425 90.585 141.205 ;
        RECT 92.275 141.035 92.445 141.725 ;
        RECT 90.945 140.865 92.445 141.035 ;
        RECT 92.635 141.065 92.845 141.855 ;
        RECT 93.015 141.235 93.365 141.855 ;
        RECT 93.535 141.245 93.705 142.025 ;
        RECT 94.235 141.865 94.405 142.095 ;
        RECT 93.875 141.695 94.405 141.865 ;
        RECT 93.875 141.415 94.095 141.695 ;
        RECT 94.575 141.525 94.815 141.925 ;
        RECT 93.535 141.075 93.940 141.245 ;
        RECT 94.275 141.155 94.815 141.525 ;
        RECT 94.985 141.740 95.305 142.095 ;
        RECT 95.550 142.015 95.855 142.475 ;
        RECT 96.025 141.765 96.280 142.295 ;
        RECT 96.455 141.930 101.800 142.475 ;
        RECT 101.975 141.930 107.320 142.475 ;
        RECT 94.985 141.565 95.310 141.740 ;
        RECT 94.985 141.265 95.900 141.565 ;
        RECT 95.160 141.235 95.900 141.265 ;
        RECT 92.635 140.905 93.310 141.065 ;
        RECT 93.770 140.985 93.940 141.075 ;
        RECT 92.635 140.895 93.600 140.905 ;
        RECT 92.275 140.725 92.445 140.865 ;
        RECT 89.020 139.925 89.270 140.385 ;
        RECT 89.440 140.095 89.690 140.425 ;
        RECT 89.905 140.095 90.585 140.425 ;
        RECT 90.755 140.525 91.830 140.695 ;
        RECT 92.275 140.555 92.835 140.725 ;
        RECT 93.140 140.605 93.600 140.895 ;
        RECT 93.770 140.815 94.990 140.985 ;
        RECT 90.755 140.185 90.925 140.525 ;
        RECT 91.160 139.925 91.490 140.355 ;
        RECT 91.660 140.185 91.830 140.525 ;
        RECT 92.125 139.925 92.495 140.385 ;
        RECT 92.665 140.095 92.835 140.555 ;
        RECT 93.770 140.435 93.940 140.815 ;
        RECT 95.160 140.645 95.330 141.235 ;
        RECT 96.070 141.115 96.280 141.765 ;
        RECT 93.070 140.095 93.940 140.435 ;
        RECT 94.530 140.475 95.330 140.645 ;
        RECT 94.110 139.925 94.360 140.385 ;
        RECT 94.530 140.185 94.700 140.475 ;
        RECT 94.880 139.925 95.210 140.305 ;
        RECT 95.550 139.925 95.855 141.065 ;
        RECT 96.025 140.235 96.280 141.115 ;
        RECT 98.040 141.100 98.380 141.930 ;
        RECT 99.860 140.360 100.210 141.610 ;
        RECT 103.560 141.100 103.900 141.930 ;
        RECT 107.955 141.725 109.165 142.475 ;
        RECT 105.380 140.360 105.730 141.610 ;
        RECT 107.955 141.015 108.475 141.555 ;
        RECT 108.645 141.185 109.165 141.725 ;
        RECT 96.455 139.925 101.800 140.360 ;
        RECT 101.975 139.925 107.320 140.360 ;
        RECT 107.955 139.925 109.165 141.015 ;
        RECT 35.190 139.755 109.250 139.925 ;
        RECT 35.275 138.665 36.485 139.755 ;
        RECT 36.655 139.320 42.000 139.755 ;
        RECT 42.175 139.320 47.520 139.755 ;
        RECT 35.275 137.955 35.795 138.495 ;
        RECT 35.965 138.125 36.485 138.665 ;
        RECT 35.275 137.205 36.485 137.955 ;
        RECT 38.240 137.750 38.580 138.580 ;
        RECT 40.060 138.070 40.410 139.320 ;
        RECT 43.760 137.750 44.100 138.580 ;
        RECT 45.580 138.070 45.930 139.320 ;
        RECT 48.155 138.590 48.445 139.755 ;
        RECT 48.615 139.320 53.960 139.755 ;
        RECT 36.655 137.205 42.000 137.750 ;
        RECT 42.175 137.205 47.520 137.750 ;
        RECT 48.155 137.205 48.445 137.930 ;
        RECT 50.200 137.750 50.540 138.580 ;
        RECT 52.020 138.070 52.370 139.320 ;
        RECT 54.135 138.665 55.345 139.755 ;
        RECT 54.135 137.955 54.655 138.495 ;
        RECT 54.825 138.125 55.345 138.665 ;
        RECT 55.555 138.615 55.785 139.755 ;
        RECT 55.955 138.605 56.285 139.585 ;
        RECT 56.455 138.615 56.665 139.755 ;
        RECT 56.895 138.665 58.565 139.755 ;
        RECT 55.535 138.195 55.865 138.445 ;
        RECT 48.615 137.205 53.960 137.750 ;
        RECT 54.135 137.205 55.345 137.955 ;
        RECT 55.555 137.205 55.785 138.025 ;
        RECT 56.035 138.005 56.285 138.605 ;
        RECT 55.955 137.375 56.285 138.005 ;
        RECT 56.455 137.205 56.665 138.025 ;
        RECT 56.895 137.975 57.645 138.495 ;
        RECT 57.815 138.145 58.565 138.665 ;
        RECT 59.195 138.955 59.635 139.585 ;
        RECT 56.895 137.205 58.565 137.975 ;
        RECT 59.195 137.945 59.505 138.955 ;
        RECT 59.810 138.905 60.125 139.755 ;
        RECT 60.295 139.415 61.725 139.585 ;
        RECT 60.295 138.735 60.465 139.415 ;
        RECT 59.675 138.565 60.465 138.735 ;
        RECT 59.675 138.115 59.845 138.565 ;
        RECT 60.635 138.445 60.835 139.245 ;
        RECT 60.015 138.115 60.405 138.395 ;
        RECT 60.590 138.115 60.835 138.445 ;
        RECT 61.035 138.115 61.285 139.245 ;
        RECT 61.475 138.785 61.725 139.415 ;
        RECT 61.905 138.955 62.235 139.755 ;
        RECT 62.415 139.285 62.755 139.545 ;
        RECT 62.925 139.295 63.175 139.755 ;
        RECT 61.475 138.615 62.245 138.785 ;
        RECT 61.500 138.115 61.905 138.445 ;
        RECT 62.075 137.945 62.245 138.615 ;
        RECT 59.195 137.385 59.635 137.945 ;
        RECT 59.805 137.205 60.255 137.945 ;
        RECT 60.425 137.775 61.585 137.945 ;
        RECT 60.425 137.375 60.595 137.775 ;
        RECT 60.765 137.205 61.185 137.605 ;
        RECT 61.355 137.375 61.585 137.775 ;
        RECT 61.755 137.375 62.245 137.945 ;
        RECT 62.415 137.680 62.675 139.285 ;
        RECT 63.365 139.115 63.695 139.545 ;
        RECT 62.845 138.945 63.695 139.115 ;
        RECT 63.865 139.085 64.035 139.585 ;
        RECT 64.245 139.295 64.495 139.755 ;
        RECT 64.705 139.085 64.875 139.585 ;
        RECT 65.175 139.295 65.425 139.755 ;
        RECT 65.665 139.085 65.835 139.585 ;
        RECT 62.845 138.025 63.015 138.945 ;
        RECT 63.865 138.915 65.835 139.085 ;
        RECT 63.335 138.195 63.665 138.755 ;
        RECT 63.865 138.445 64.165 138.740 ;
        RECT 63.865 138.395 64.245 138.445 ;
        RECT 63.855 138.225 64.245 138.395 ;
        RECT 63.865 138.115 64.245 138.225 ;
        RECT 62.845 137.930 63.665 138.025 ;
        RECT 62.845 137.855 63.860 137.930 ;
        RECT 62.415 137.420 62.755 137.680 ;
        RECT 62.925 137.205 63.255 137.685 ;
        RECT 63.445 137.420 63.860 137.855 ;
        RECT 64.555 137.720 64.775 138.445 ;
        RECT 65.035 138.115 65.415 138.745 ;
        RECT 65.645 138.115 65.900 138.745 ;
        RECT 66.095 138.615 66.480 139.585 ;
        RECT 66.650 139.295 66.975 139.755 ;
        RECT 67.495 139.125 67.775 139.585 ;
        RECT 66.650 138.905 67.775 139.125 ;
        RECT 64.030 137.535 64.980 137.720 ;
        RECT 65.210 137.515 65.415 138.115 ;
        RECT 66.095 137.945 66.375 138.615 ;
        RECT 66.650 138.445 67.100 138.905 ;
        RECT 67.965 138.735 68.365 139.585 ;
        RECT 68.765 139.295 69.035 139.755 ;
        RECT 69.205 139.125 69.490 139.585 ;
        RECT 70.275 139.295 70.490 139.755 ;
        RECT 70.660 139.125 70.990 139.585 ;
        RECT 66.545 138.115 67.100 138.445 ;
        RECT 67.270 138.175 68.365 138.735 ;
        RECT 66.650 138.005 67.100 138.115 ;
        RECT 65.585 137.205 65.925 137.930 ;
        RECT 66.095 137.375 66.480 137.945 ;
        RECT 66.650 137.835 67.775 138.005 ;
        RECT 66.650 137.205 66.975 137.665 ;
        RECT 67.495 137.375 67.775 137.835 ;
        RECT 67.965 137.375 68.365 138.175 ;
        RECT 68.535 138.905 69.490 139.125 ;
        RECT 69.820 138.955 70.990 139.125 ;
        RECT 71.160 138.955 71.410 139.755 ;
        RECT 68.535 138.005 68.745 138.905 ;
        RECT 68.915 138.175 69.605 138.735 ;
        RECT 68.535 137.835 69.490 138.005 ;
        RECT 68.765 137.205 69.035 137.665 ;
        RECT 69.205 137.375 69.490 137.835 ;
        RECT 69.820 137.665 70.190 138.955 ;
        RECT 71.620 138.785 71.900 138.945 ;
        RECT 70.565 138.615 71.900 138.785 ;
        RECT 72.075 138.665 73.745 139.755 ;
        RECT 70.565 138.445 70.735 138.615 ;
        RECT 70.360 138.195 70.735 138.445 ;
        RECT 70.905 138.195 71.380 138.435 ;
        RECT 71.550 138.195 71.900 138.435 ;
        RECT 70.565 138.025 70.735 138.195 ;
        RECT 70.565 137.855 71.900 138.025 ;
        RECT 69.820 137.375 70.570 137.665 ;
        RECT 71.080 137.205 71.410 137.665 ;
        RECT 71.630 137.645 71.900 137.855 ;
        RECT 72.075 137.975 72.825 138.495 ;
        RECT 72.995 138.145 73.745 138.665 ;
        RECT 73.915 138.590 74.205 139.755 ;
        RECT 74.375 138.665 75.585 139.755 ;
        RECT 72.075 137.205 73.745 137.975 ;
        RECT 74.375 137.955 74.895 138.495 ;
        RECT 75.065 138.125 75.585 138.665 ;
        RECT 75.765 138.615 76.095 139.755 ;
        RECT 76.625 138.785 76.955 139.570 ;
        RECT 76.275 138.615 76.955 138.785 ;
        RECT 77.160 138.785 77.460 138.980 ;
        RECT 77.630 138.955 77.885 139.755 ;
        RECT 78.085 139.125 78.415 139.585 ;
        RECT 78.585 139.295 79.160 139.755 ;
        RECT 79.330 139.125 79.685 139.585 ;
        RECT 78.085 138.955 79.685 139.125 ;
        RECT 77.160 138.615 78.410 138.785 ;
        RECT 75.755 138.195 76.105 138.445 ;
        RECT 76.275 138.015 76.445 138.615 ;
        RECT 76.615 138.195 76.965 138.445 ;
        RECT 73.915 137.205 74.205 137.930 ;
        RECT 74.375 137.205 75.585 137.955 ;
        RECT 75.765 137.205 76.035 138.015 ;
        RECT 76.205 137.375 76.535 138.015 ;
        RECT 76.705 137.205 76.945 138.015 ;
        RECT 77.160 137.960 77.330 138.615 ;
        RECT 77.505 138.115 77.850 138.445 ;
        RECT 78.080 138.195 78.410 138.615 ;
        RECT 78.580 138.025 78.860 138.955 ;
        RECT 79.040 138.395 79.230 138.775 ;
        RECT 79.410 138.615 79.685 138.955 ;
        RECT 79.855 138.615 80.185 139.755 ;
        RECT 80.365 138.945 80.660 139.755 ;
        RECT 80.840 138.445 81.085 139.585 ;
        RECT 81.260 138.945 81.520 139.755 ;
        RECT 82.120 139.750 88.395 139.755 ;
        RECT 81.700 138.445 81.950 139.580 ;
        RECT 82.120 138.955 82.380 139.750 ;
        RECT 82.550 138.855 82.810 139.580 ;
        RECT 82.980 139.025 83.240 139.750 ;
        RECT 83.410 138.855 83.670 139.580 ;
        RECT 83.840 139.025 84.100 139.750 ;
        RECT 84.270 138.855 84.530 139.580 ;
        RECT 84.700 139.025 84.960 139.750 ;
        RECT 85.130 138.855 85.390 139.580 ;
        RECT 85.560 139.025 85.805 139.750 ;
        RECT 85.975 138.855 86.235 139.580 ;
        RECT 86.420 139.025 86.665 139.750 ;
        RECT 86.835 138.855 87.095 139.580 ;
        RECT 87.280 139.025 87.525 139.750 ;
        RECT 87.695 138.855 87.955 139.580 ;
        RECT 88.140 139.025 88.395 139.750 ;
        RECT 82.550 138.840 87.955 138.855 ;
        RECT 88.565 138.840 88.855 139.580 ;
        RECT 89.025 139.010 89.295 139.755 ;
        RECT 82.550 138.615 89.295 138.840 ;
        RECT 79.035 138.225 80.185 138.395 ;
        RECT 79.040 138.195 80.185 138.225 ;
        RECT 77.160 137.630 77.395 137.960 ;
        RECT 77.565 137.205 77.895 137.945 ;
        RECT 78.130 137.585 78.405 138.025 ;
        RECT 78.580 137.925 78.905 138.025 ;
        RECT 78.575 137.755 78.905 137.925 ;
        RECT 79.075 137.815 80.185 138.025 ;
        RECT 80.355 137.885 80.670 138.445 ;
        RECT 80.840 138.195 87.960 138.445 ;
        RECT 79.075 137.585 79.325 137.815 ;
        RECT 78.130 137.375 79.325 137.585 ;
        RECT 79.495 137.205 79.665 137.645 ;
        RECT 79.835 137.375 80.185 137.815 ;
        RECT 80.355 137.205 80.660 137.715 ;
        RECT 80.840 137.385 81.090 138.195 ;
        RECT 81.260 137.205 81.520 137.730 ;
        RECT 81.700 137.385 81.950 138.195 ;
        RECT 88.130 138.025 89.295 138.615 ;
        RECT 82.550 137.855 89.295 138.025 ;
        RECT 89.555 138.615 89.940 139.585 ;
        RECT 90.110 139.295 90.435 139.755 ;
        RECT 90.955 139.125 91.235 139.585 ;
        RECT 90.110 138.905 91.235 139.125 ;
        RECT 89.555 137.945 89.835 138.615 ;
        RECT 90.110 138.445 90.560 138.905 ;
        RECT 91.425 138.735 91.825 139.585 ;
        RECT 92.225 139.295 92.495 139.755 ;
        RECT 92.665 139.125 92.950 139.585 ;
        RECT 90.005 138.115 90.560 138.445 ;
        RECT 90.730 138.175 91.825 138.735 ;
        RECT 90.110 138.005 90.560 138.115 ;
        RECT 82.120 137.205 82.380 137.765 ;
        RECT 82.550 137.400 82.810 137.855 ;
        RECT 82.980 137.205 83.240 137.685 ;
        RECT 83.410 137.400 83.670 137.855 ;
        RECT 83.840 137.205 84.100 137.685 ;
        RECT 84.270 137.400 84.530 137.855 ;
        RECT 84.700 137.205 84.945 137.685 ;
        RECT 85.115 137.400 85.390 137.855 ;
        RECT 85.560 137.205 85.805 137.685 ;
        RECT 85.975 137.400 86.235 137.855 ;
        RECT 86.415 137.205 86.665 137.685 ;
        RECT 86.835 137.400 87.095 137.855 ;
        RECT 87.275 137.205 87.525 137.685 ;
        RECT 87.695 137.400 87.955 137.855 ;
        RECT 88.135 137.205 88.395 137.685 ;
        RECT 88.565 137.400 88.825 137.855 ;
        RECT 88.995 137.205 89.295 137.685 ;
        RECT 89.555 137.375 89.940 137.945 ;
        RECT 90.110 137.835 91.235 138.005 ;
        RECT 90.110 137.205 90.435 137.665 ;
        RECT 90.955 137.375 91.235 137.835 ;
        RECT 91.425 137.375 91.825 138.175 ;
        RECT 91.995 138.905 92.950 139.125 ;
        RECT 91.995 138.005 92.205 138.905 ;
        RECT 92.375 138.175 93.065 138.735 ;
        RECT 93.240 138.615 93.560 139.755 ;
        RECT 93.740 138.445 93.935 139.495 ;
        RECT 94.115 138.905 94.445 139.585 ;
        RECT 94.645 138.955 94.900 139.755 ;
        RECT 94.115 138.625 94.465 138.905 ;
        RECT 93.300 138.395 93.560 138.445 ;
        RECT 93.295 138.225 93.560 138.395 ;
        RECT 93.300 138.115 93.560 138.225 ;
        RECT 93.740 138.115 94.125 138.445 ;
        RECT 94.295 138.245 94.465 138.625 ;
        RECT 94.655 138.415 94.900 138.775 ;
        RECT 95.115 138.615 95.345 139.755 ;
        RECT 95.515 138.605 95.845 139.585 ;
        RECT 96.015 138.615 96.225 139.755 ;
        RECT 96.455 138.665 99.045 139.755 ;
        RECT 94.295 138.075 94.815 138.245 ;
        RECT 95.095 138.195 95.425 138.445 ;
        RECT 91.995 137.835 92.950 138.005 ;
        RECT 92.225 137.205 92.495 137.665 ;
        RECT 92.665 137.375 92.950 137.835 ;
        RECT 93.240 137.735 94.455 137.905 ;
        RECT 93.240 137.385 93.530 137.735 ;
        RECT 93.725 137.205 94.055 137.565 ;
        RECT 94.225 137.430 94.455 137.735 ;
        RECT 94.645 137.510 94.815 138.075 ;
        RECT 95.115 137.205 95.345 138.025 ;
        RECT 95.595 138.005 95.845 138.605 ;
        RECT 95.515 137.375 95.845 138.005 ;
        RECT 96.015 137.205 96.225 138.025 ;
        RECT 96.455 137.975 97.665 138.495 ;
        RECT 97.835 138.145 99.045 138.665 ;
        RECT 99.675 138.590 99.965 139.755 ;
        RECT 100.135 138.665 103.645 139.755 ;
        RECT 100.135 137.975 101.785 138.495 ;
        RECT 101.955 138.145 103.645 138.665 ;
        RECT 104.775 138.615 105.005 139.755 ;
        RECT 105.175 138.605 105.505 139.585 ;
        RECT 105.675 138.615 105.885 139.755 ;
        RECT 106.115 138.665 107.785 139.755 ;
        RECT 104.755 138.195 105.085 138.445 ;
        RECT 96.455 137.205 99.045 137.975 ;
        RECT 99.675 137.205 99.965 137.930 ;
        RECT 100.135 137.205 103.645 137.975 ;
        RECT 104.775 137.205 105.005 138.025 ;
        RECT 105.255 138.005 105.505 138.605 ;
        RECT 105.175 137.375 105.505 138.005 ;
        RECT 105.675 137.205 105.885 138.025 ;
        RECT 106.115 137.975 106.865 138.495 ;
        RECT 107.035 138.145 107.785 138.665 ;
        RECT 107.955 138.665 109.165 139.755 ;
        RECT 107.955 138.125 108.475 138.665 ;
        RECT 106.115 137.205 107.785 137.975 ;
        RECT 108.645 137.955 109.165 138.495 ;
        RECT 107.955 137.205 109.165 137.955 ;
        RECT 35.190 137.035 109.250 137.205 ;
        RECT 35.275 136.285 36.485 137.035 ;
        RECT 36.655 136.490 42.000 137.035 ;
        RECT 42.175 136.490 47.520 137.035 ;
        RECT 35.275 135.745 35.795 136.285 ;
        RECT 35.965 135.575 36.485 136.115 ;
        RECT 38.240 135.660 38.580 136.490 ;
        RECT 35.275 134.485 36.485 135.575 ;
        RECT 40.060 134.920 40.410 136.170 ;
        RECT 43.760 135.660 44.100 136.490 ;
        RECT 47.695 136.265 51.205 137.035 ;
        RECT 51.840 136.485 52.095 136.775 ;
        RECT 52.265 136.655 52.595 137.035 ;
        RECT 51.840 136.315 52.590 136.485 ;
        RECT 45.580 134.920 45.930 136.170 ;
        RECT 47.695 135.745 49.345 136.265 ;
        RECT 49.515 135.575 51.205 136.095 ;
        RECT 36.655 134.485 42.000 134.920 ;
        RECT 42.175 134.485 47.520 134.920 ;
        RECT 47.695 134.485 51.205 135.575 ;
        RECT 51.840 135.495 52.190 136.145 ;
        RECT 52.360 135.325 52.590 136.315 ;
        RECT 51.840 135.155 52.590 135.325 ;
        RECT 51.840 134.655 52.095 135.155 ;
        RECT 52.265 134.485 52.595 134.985 ;
        RECT 52.765 134.655 52.935 136.775 ;
        RECT 53.295 136.675 53.625 137.035 ;
        RECT 53.795 136.645 54.290 136.815 ;
        RECT 54.495 136.645 55.350 136.815 ;
        RECT 53.165 135.455 53.625 136.505 ;
        RECT 53.105 134.670 53.430 135.455 ;
        RECT 53.795 135.285 53.965 136.645 ;
        RECT 54.135 135.735 54.485 136.355 ;
        RECT 54.655 136.135 55.010 136.355 ;
        RECT 54.655 135.545 54.825 136.135 ;
        RECT 55.180 135.935 55.350 136.645 ;
        RECT 56.225 136.575 56.555 137.035 ;
        RECT 56.765 136.675 57.115 136.845 ;
        RECT 55.555 136.105 56.345 136.355 ;
        RECT 56.765 136.285 57.025 136.675 ;
        RECT 57.335 136.585 58.285 136.865 ;
        RECT 58.455 136.595 58.645 137.035 ;
        RECT 58.815 136.655 59.885 136.825 ;
        RECT 56.515 135.935 56.685 136.115 ;
        RECT 53.795 135.115 54.190 135.285 ;
        RECT 54.360 135.155 54.825 135.545 ;
        RECT 54.995 135.765 56.685 135.935 ;
        RECT 54.020 134.985 54.190 135.115 ;
        RECT 54.995 134.985 55.165 135.765 ;
        RECT 56.855 135.595 57.025 136.285 ;
        RECT 55.525 135.425 57.025 135.595 ;
        RECT 57.215 135.625 57.425 136.415 ;
        RECT 57.595 135.795 57.945 136.415 ;
        RECT 58.115 135.805 58.285 136.585 ;
        RECT 58.815 136.425 58.985 136.655 ;
        RECT 58.455 136.255 58.985 136.425 ;
        RECT 58.455 135.975 58.675 136.255 ;
        RECT 59.155 136.085 59.395 136.485 ;
        RECT 58.115 135.635 58.520 135.805 ;
        RECT 58.855 135.715 59.395 136.085 ;
        RECT 59.565 136.300 59.885 136.655 ;
        RECT 60.130 136.575 60.435 137.035 ;
        RECT 60.605 136.325 60.860 136.855 ;
        RECT 59.565 136.125 59.890 136.300 ;
        RECT 59.565 135.825 60.480 136.125 ;
        RECT 59.740 135.795 60.480 135.825 ;
        RECT 57.215 135.465 57.890 135.625 ;
        RECT 58.350 135.545 58.520 135.635 ;
        RECT 57.215 135.455 58.180 135.465 ;
        RECT 56.855 135.285 57.025 135.425 ;
        RECT 53.600 134.485 53.850 134.945 ;
        RECT 54.020 134.655 54.270 134.985 ;
        RECT 54.485 134.655 55.165 134.985 ;
        RECT 55.335 135.085 56.410 135.255 ;
        RECT 56.855 135.115 57.415 135.285 ;
        RECT 57.720 135.165 58.180 135.455 ;
        RECT 58.350 135.375 59.570 135.545 ;
        RECT 55.335 134.745 55.505 135.085 ;
        RECT 55.740 134.485 56.070 134.915 ;
        RECT 56.240 134.745 56.410 135.085 ;
        RECT 56.705 134.485 57.075 134.945 ;
        RECT 57.245 134.655 57.415 135.115 ;
        RECT 58.350 134.995 58.520 135.375 ;
        RECT 59.740 135.205 59.910 135.795 ;
        RECT 60.650 135.675 60.860 136.325 ;
        RECT 61.035 136.310 61.325 137.035 ;
        RECT 61.555 136.215 61.765 137.035 ;
        RECT 61.935 136.235 62.265 136.865 ;
        RECT 57.650 134.655 58.520 134.995 ;
        RECT 59.110 135.035 59.910 135.205 ;
        RECT 58.690 134.485 58.940 134.945 ;
        RECT 59.110 134.745 59.280 135.035 ;
        RECT 59.460 134.485 59.790 134.865 ;
        RECT 60.130 134.485 60.435 135.625 ;
        RECT 60.605 134.795 60.860 135.675 ;
        RECT 61.035 134.485 61.325 135.650 ;
        RECT 61.935 135.635 62.185 136.235 ;
        RECT 62.435 136.215 62.665 137.035 ;
        RECT 62.875 136.265 65.465 137.035 ;
        RECT 62.355 135.795 62.685 136.045 ;
        RECT 62.875 135.745 64.085 136.265 ;
        RECT 66.135 136.215 66.365 137.035 ;
        RECT 66.535 136.235 66.865 136.865 ;
        RECT 61.555 134.485 61.765 135.625 ;
        RECT 61.935 134.655 62.265 135.635 ;
        RECT 62.435 134.485 62.665 135.625 ;
        RECT 64.255 135.575 65.465 136.095 ;
        RECT 66.115 135.795 66.445 136.045 ;
        RECT 66.615 135.635 66.865 136.235 ;
        RECT 67.035 136.215 67.245 137.035 ;
        RECT 67.475 136.265 70.065 137.035 ;
        RECT 70.350 136.405 70.635 136.865 ;
        RECT 70.805 136.575 71.075 137.035 ;
        RECT 67.475 135.745 68.685 136.265 ;
        RECT 70.350 136.235 71.305 136.405 ;
        RECT 62.875 134.485 65.465 135.575 ;
        RECT 66.135 134.485 66.365 135.625 ;
        RECT 66.535 134.655 66.865 135.635 ;
        RECT 67.035 134.485 67.245 135.625 ;
        RECT 68.855 135.575 70.065 136.095 ;
        RECT 67.475 134.485 70.065 135.575 ;
        RECT 70.235 135.505 70.925 136.065 ;
        RECT 71.095 135.335 71.305 136.235 ;
        RECT 70.350 135.115 71.305 135.335 ;
        RECT 71.475 136.065 71.875 136.865 ;
        RECT 72.065 136.405 72.345 136.865 ;
        RECT 72.865 136.575 73.190 137.035 ;
        RECT 72.065 136.235 73.190 136.405 ;
        RECT 73.360 136.295 73.745 136.865 ;
        RECT 73.935 136.305 74.225 137.035 ;
        RECT 72.740 136.125 73.190 136.235 ;
        RECT 71.475 135.505 72.570 136.065 ;
        RECT 72.740 135.795 73.295 136.125 ;
        RECT 70.350 134.655 70.635 135.115 ;
        RECT 70.805 134.485 71.075 134.945 ;
        RECT 71.475 134.655 71.875 135.505 ;
        RECT 72.740 135.335 73.190 135.795 ;
        RECT 73.465 135.625 73.745 136.295 ;
        RECT 73.925 135.795 74.225 136.125 ;
        RECT 74.405 136.105 74.635 136.745 ;
        RECT 74.815 136.485 75.125 136.855 ;
        RECT 75.305 136.665 75.975 137.035 ;
        RECT 74.815 136.285 76.045 136.485 ;
        RECT 74.405 135.795 74.930 136.105 ;
        RECT 75.110 135.795 75.575 136.105 ;
        RECT 72.065 135.115 73.190 135.335 ;
        RECT 72.065 134.655 72.345 135.115 ;
        RECT 72.865 134.485 73.190 134.945 ;
        RECT 73.360 134.655 73.745 135.625 ;
        RECT 75.755 135.615 76.045 136.285 ;
        RECT 73.935 135.375 75.095 135.615 ;
        RECT 73.935 134.665 74.195 135.375 ;
        RECT 74.365 134.485 74.695 135.195 ;
        RECT 74.865 134.665 75.095 135.375 ;
        RECT 75.275 135.395 76.045 135.615 ;
        RECT 75.275 134.665 75.545 135.395 ;
        RECT 75.725 134.485 76.065 135.215 ;
        RECT 76.235 134.665 76.495 136.855 ;
        RECT 77.600 136.505 77.890 136.855 ;
        RECT 78.085 136.675 78.415 137.035 ;
        RECT 78.585 136.505 78.815 136.810 ;
        RECT 77.600 136.335 78.815 136.505 ;
        RECT 79.005 136.165 79.175 136.730 ;
        RECT 79.445 136.535 79.775 137.035 ;
        RECT 79.975 136.465 80.145 136.815 ;
        RECT 80.345 136.635 80.675 137.035 ;
        RECT 80.845 136.465 81.015 136.815 ;
        RECT 81.185 136.635 81.565 137.035 ;
        RECT 77.660 136.015 77.920 136.125 ;
        RECT 77.655 135.845 77.920 136.015 ;
        RECT 77.660 135.795 77.920 135.845 ;
        RECT 78.100 135.795 78.485 136.125 ;
        RECT 78.655 135.995 79.175 136.165 ;
        RECT 77.600 134.485 77.920 135.625 ;
        RECT 78.100 134.745 78.295 135.795 ;
        RECT 78.655 135.615 78.825 135.995 ;
        RECT 78.475 135.335 78.825 135.615 ;
        RECT 79.015 135.465 79.260 135.825 ;
        RECT 79.440 135.795 79.790 136.365 ;
        RECT 79.975 136.295 81.585 136.465 ;
        RECT 81.755 136.360 82.025 136.705 ;
        RECT 81.415 136.125 81.585 136.295 ;
        RECT 79.440 135.335 79.760 135.625 ;
        RECT 79.960 135.505 80.670 136.125 ;
        RECT 80.840 135.795 81.245 136.125 ;
        RECT 81.415 135.795 81.685 136.125 ;
        RECT 81.415 135.625 81.585 135.795 ;
        RECT 81.855 135.625 82.025 136.360 ;
        RECT 82.205 136.315 82.535 137.035 ;
        RECT 83.080 136.635 84.695 136.805 ;
        RECT 84.865 136.635 85.195 137.035 ;
        RECT 84.525 136.465 84.695 136.635 ;
        RECT 85.365 136.560 85.700 136.820 ;
        RECT 82.260 136.015 82.610 136.125 ;
        RECT 82.255 135.845 82.610 136.015 ;
        RECT 80.860 135.455 81.585 135.625 ;
        RECT 80.860 135.335 81.030 135.455 ;
        RECT 78.475 134.655 78.805 135.335 ;
        RECT 79.005 134.485 79.260 135.285 ;
        RECT 79.440 135.165 81.030 135.335 ;
        RECT 79.440 134.705 81.095 134.995 ;
        RECT 81.265 134.485 81.545 135.285 ;
        RECT 81.755 134.655 82.025 135.625 ;
        RECT 82.260 135.795 82.610 135.845 ;
        RECT 82.920 135.795 83.340 136.460 ;
        RECT 83.510 136.015 83.800 136.455 ;
        RECT 83.990 136.355 84.260 136.455 ;
        RECT 83.990 136.185 84.265 136.355 ;
        RECT 84.525 136.295 85.085 136.465 ;
        RECT 83.510 135.845 83.805 136.015 ;
        RECT 83.510 135.795 83.800 135.845 ;
        RECT 83.990 135.795 84.260 136.185 ;
        RECT 84.915 136.125 85.085 136.295 ;
        RECT 84.470 136.015 84.720 136.125 ;
        RECT 84.470 135.845 84.725 136.015 ;
        RECT 84.470 135.795 84.720 135.845 ;
        RECT 84.915 135.795 85.220 136.125 ;
        RECT 82.260 135.505 82.465 135.795 ;
        RECT 84.915 135.625 85.085 135.795 ;
        RECT 82.715 135.455 85.085 135.625 ;
        RECT 82.285 134.825 82.455 135.325 ;
        RECT 82.715 134.995 82.885 135.455 ;
        RECT 83.115 135.075 84.540 135.245 ;
        RECT 83.115 134.825 83.445 135.075 ;
        RECT 82.285 134.655 83.445 134.825 ;
        RECT 83.670 134.485 84.000 134.905 ;
        RECT 84.255 134.655 84.540 135.075 ;
        RECT 84.785 134.485 85.115 135.285 ;
        RECT 85.445 135.205 85.700 136.560 ;
        RECT 86.795 136.310 87.085 137.035 ;
        RECT 87.260 136.485 87.515 136.775 ;
        RECT 87.685 136.655 88.015 137.035 ;
        RECT 87.260 136.315 88.010 136.485 ;
        RECT 85.365 134.695 85.700 135.205 ;
        RECT 86.795 134.485 87.085 135.650 ;
        RECT 87.260 135.495 87.610 136.145 ;
        RECT 87.780 135.325 88.010 136.315 ;
        RECT 87.260 135.155 88.010 135.325 ;
        RECT 87.260 134.655 87.515 135.155 ;
        RECT 87.685 134.485 88.015 134.985 ;
        RECT 88.185 134.655 88.355 136.775 ;
        RECT 88.715 136.675 89.045 137.035 ;
        RECT 89.215 136.645 89.710 136.815 ;
        RECT 89.915 136.645 90.770 136.815 ;
        RECT 88.585 135.455 89.045 136.505 ;
        RECT 88.525 134.670 88.850 135.455 ;
        RECT 89.215 135.285 89.385 136.645 ;
        RECT 89.555 135.735 89.905 136.355 ;
        RECT 90.075 136.135 90.430 136.355 ;
        RECT 90.075 135.545 90.245 136.135 ;
        RECT 90.600 135.935 90.770 136.645 ;
        RECT 91.645 136.575 91.975 137.035 ;
        RECT 92.185 136.675 92.535 136.845 ;
        RECT 90.975 136.105 91.765 136.355 ;
        RECT 92.185 136.285 92.445 136.675 ;
        RECT 92.755 136.585 93.705 136.865 ;
        RECT 93.875 136.595 94.065 137.035 ;
        RECT 94.235 136.655 95.305 136.825 ;
        RECT 91.935 135.935 92.105 136.115 ;
        RECT 89.215 135.115 89.610 135.285 ;
        RECT 89.780 135.155 90.245 135.545 ;
        RECT 90.415 135.765 92.105 135.935 ;
        RECT 89.440 134.985 89.610 135.115 ;
        RECT 90.415 134.985 90.585 135.765 ;
        RECT 92.275 135.595 92.445 136.285 ;
        RECT 90.945 135.425 92.445 135.595 ;
        RECT 92.635 135.625 92.845 136.415 ;
        RECT 93.015 135.795 93.365 136.415 ;
        RECT 93.535 135.805 93.705 136.585 ;
        RECT 94.235 136.425 94.405 136.655 ;
        RECT 93.875 136.255 94.405 136.425 ;
        RECT 93.875 135.975 94.095 136.255 ;
        RECT 94.575 136.085 94.815 136.485 ;
        RECT 93.535 135.635 93.940 135.805 ;
        RECT 94.275 135.715 94.815 136.085 ;
        RECT 94.985 136.300 95.305 136.655 ;
        RECT 95.550 136.575 95.855 137.035 ;
        RECT 96.025 136.325 96.280 136.855 ;
        RECT 96.455 136.490 101.800 137.035 ;
        RECT 101.975 136.490 107.320 137.035 ;
        RECT 94.985 136.125 95.310 136.300 ;
        RECT 94.985 135.825 95.900 136.125 ;
        RECT 95.160 135.795 95.900 135.825 ;
        RECT 92.635 135.465 93.310 135.625 ;
        RECT 93.770 135.545 93.940 135.635 ;
        RECT 92.635 135.455 93.600 135.465 ;
        RECT 92.275 135.285 92.445 135.425 ;
        RECT 89.020 134.485 89.270 134.945 ;
        RECT 89.440 134.655 89.690 134.985 ;
        RECT 89.905 134.655 90.585 134.985 ;
        RECT 90.755 135.085 91.830 135.255 ;
        RECT 92.275 135.115 92.835 135.285 ;
        RECT 93.140 135.165 93.600 135.455 ;
        RECT 93.770 135.375 94.990 135.545 ;
        RECT 90.755 134.745 90.925 135.085 ;
        RECT 91.160 134.485 91.490 134.915 ;
        RECT 91.660 134.745 91.830 135.085 ;
        RECT 92.125 134.485 92.495 134.945 ;
        RECT 92.665 134.655 92.835 135.115 ;
        RECT 93.770 134.995 93.940 135.375 ;
        RECT 95.160 135.205 95.330 135.795 ;
        RECT 96.070 135.675 96.280 136.325 ;
        RECT 93.070 134.655 93.940 134.995 ;
        RECT 94.530 135.035 95.330 135.205 ;
        RECT 94.110 134.485 94.360 134.945 ;
        RECT 94.530 134.745 94.700 135.035 ;
        RECT 94.880 134.485 95.210 134.865 ;
        RECT 95.550 134.485 95.855 135.625 ;
        RECT 96.025 134.795 96.280 135.675 ;
        RECT 98.040 135.660 98.380 136.490 ;
        RECT 99.860 134.920 100.210 136.170 ;
        RECT 103.560 135.660 103.900 136.490 ;
        RECT 107.955 136.285 109.165 137.035 ;
        RECT 105.380 134.920 105.730 136.170 ;
        RECT 107.955 135.575 108.475 136.115 ;
        RECT 108.645 135.745 109.165 136.285 ;
        RECT 96.455 134.485 101.800 134.920 ;
        RECT 101.975 134.485 107.320 134.920 ;
        RECT 107.955 134.485 109.165 135.575 ;
        RECT 35.190 134.315 109.250 134.485 ;
        RECT 35.275 133.225 36.485 134.315 ;
        RECT 36.655 133.880 42.000 134.315 ;
        RECT 42.175 133.880 47.520 134.315 ;
        RECT 35.275 132.515 35.795 133.055 ;
        RECT 35.965 132.685 36.485 133.225 ;
        RECT 35.275 131.765 36.485 132.515 ;
        RECT 38.240 132.310 38.580 133.140 ;
        RECT 40.060 132.630 40.410 133.880 ;
        RECT 43.760 132.310 44.100 133.140 ;
        RECT 45.580 132.630 45.930 133.880 ;
        RECT 48.155 133.150 48.445 134.315 ;
        RECT 48.615 133.880 53.960 134.315 ;
        RECT 54.135 133.880 59.480 134.315 ;
        RECT 36.655 131.765 42.000 132.310 ;
        RECT 42.175 131.765 47.520 132.310 ;
        RECT 48.155 131.765 48.445 132.490 ;
        RECT 50.200 132.310 50.540 133.140 ;
        RECT 52.020 132.630 52.370 133.880 ;
        RECT 55.720 132.310 56.060 133.140 ;
        RECT 57.540 132.630 57.890 133.880 ;
        RECT 59.655 133.225 61.325 134.315 ;
        RECT 61.585 133.645 61.755 134.145 ;
        RECT 61.925 133.815 62.255 134.315 ;
        RECT 61.585 133.475 62.250 133.645 ;
        RECT 59.655 132.535 60.405 133.055 ;
        RECT 60.575 132.705 61.325 133.225 ;
        RECT 61.500 132.655 61.850 133.305 ;
        RECT 48.615 131.765 53.960 132.310 ;
        RECT 54.135 131.765 59.480 132.310 ;
        RECT 59.655 131.765 61.325 132.535 ;
        RECT 62.020 132.485 62.250 133.475 ;
        RECT 61.585 132.315 62.250 132.485 ;
        RECT 61.585 132.025 61.755 132.315 ;
        RECT 61.925 131.765 62.255 132.145 ;
        RECT 62.425 132.025 62.650 134.145 ;
        RECT 62.865 133.815 63.195 134.315 ;
        RECT 63.365 133.645 63.535 134.145 ;
        RECT 63.770 133.930 64.600 134.100 ;
        RECT 64.840 133.935 65.220 134.315 ;
        RECT 62.840 133.475 63.535 133.645 ;
        RECT 62.840 132.505 63.010 133.475 ;
        RECT 63.180 132.685 63.590 133.305 ;
        RECT 63.760 133.255 64.260 133.635 ;
        RECT 62.840 132.315 63.535 132.505 ;
        RECT 63.760 132.385 63.980 133.255 ;
        RECT 64.430 133.085 64.600 133.930 ;
        RECT 65.400 133.765 65.570 134.055 ;
        RECT 65.740 133.935 66.070 134.315 ;
        RECT 66.540 133.845 67.170 134.095 ;
        RECT 67.350 133.935 67.770 134.315 ;
        RECT 67.000 133.765 67.170 133.845 ;
        RECT 67.970 133.765 68.210 134.055 ;
        RECT 64.770 133.515 66.140 133.765 ;
        RECT 64.770 133.255 65.020 133.515 ;
        RECT 65.530 133.085 65.780 133.245 ;
        RECT 64.430 132.915 65.780 133.085 ;
        RECT 64.430 132.875 64.850 132.915 ;
        RECT 64.160 132.325 64.510 132.695 ;
        RECT 62.865 131.765 63.195 132.145 ;
        RECT 63.365 131.985 63.535 132.315 ;
        RECT 64.680 132.145 64.850 132.875 ;
        RECT 65.950 132.745 66.140 133.515 ;
        RECT 65.020 132.415 65.430 132.745 ;
        RECT 65.720 132.405 66.140 132.745 ;
        RECT 66.310 133.335 66.830 133.645 ;
        RECT 67.000 133.595 68.210 133.765 ;
        RECT 68.440 133.625 68.770 134.315 ;
        RECT 66.310 132.575 66.480 133.335 ;
        RECT 66.650 132.745 66.830 133.155 ;
        RECT 67.000 133.085 67.170 133.595 ;
        RECT 68.940 133.445 69.110 134.055 ;
        RECT 69.380 133.595 69.710 134.105 ;
        RECT 68.940 133.425 69.260 133.445 ;
        RECT 67.340 133.255 69.260 133.425 ;
        RECT 67.000 132.915 68.900 133.085 ;
        RECT 67.230 132.575 67.560 132.695 ;
        RECT 66.310 132.405 67.560 132.575 ;
        RECT 63.835 131.945 64.850 132.145 ;
        RECT 65.020 131.765 65.430 132.205 ;
        RECT 65.720 131.975 65.970 132.405 ;
        RECT 66.170 131.765 66.490 132.225 ;
        RECT 67.730 132.155 67.900 132.915 ;
        RECT 68.570 132.855 68.900 132.915 ;
        RECT 68.090 132.685 68.420 132.745 ;
        RECT 68.090 132.415 68.750 132.685 ;
        RECT 69.070 132.360 69.260 133.255 ;
        RECT 67.050 131.985 67.900 132.155 ;
        RECT 68.100 131.765 68.760 132.245 ;
        RECT 68.940 132.030 69.260 132.360 ;
        RECT 69.460 133.005 69.710 133.595 ;
        RECT 69.890 133.515 70.175 134.315 ;
        RECT 70.355 133.335 70.610 134.005 ;
        RECT 70.430 133.295 70.610 133.335 ;
        RECT 70.430 133.125 70.695 133.295 ;
        RECT 71.155 133.225 72.365 134.315 ;
        RECT 69.460 132.675 70.260 133.005 ;
        RECT 69.460 132.025 69.710 132.675 ;
        RECT 70.430 132.475 70.610 133.125 ;
        RECT 69.890 131.765 70.175 132.225 ;
        RECT 70.355 131.945 70.610 132.475 ;
        RECT 71.155 132.515 71.675 133.055 ;
        RECT 71.845 132.685 72.365 133.225 ;
        RECT 72.595 133.175 72.805 134.315 ;
        RECT 72.975 133.165 73.305 134.145 ;
        RECT 73.475 133.175 73.705 134.315 ;
        RECT 71.155 131.765 72.365 132.515 ;
        RECT 72.595 131.765 72.805 132.585 ;
        RECT 72.975 132.565 73.225 133.165 ;
        RECT 73.915 133.150 74.205 134.315 ;
        RECT 74.375 133.175 74.760 134.145 ;
        RECT 74.930 133.855 75.255 134.315 ;
        RECT 75.775 133.685 76.055 134.145 ;
        RECT 74.930 133.465 76.055 133.685 ;
        RECT 73.395 132.755 73.725 133.005 ;
        RECT 72.975 131.935 73.305 132.565 ;
        RECT 73.475 131.765 73.705 132.585 ;
        RECT 74.375 132.505 74.655 133.175 ;
        RECT 74.930 133.005 75.380 133.465 ;
        RECT 76.245 133.295 76.645 134.145 ;
        RECT 77.045 133.855 77.315 134.315 ;
        RECT 77.485 133.685 77.770 134.145 ;
        RECT 74.825 132.675 75.380 133.005 ;
        RECT 75.550 132.735 76.645 133.295 ;
        RECT 74.930 132.565 75.380 132.675 ;
        RECT 73.915 131.765 74.205 132.490 ;
        RECT 74.375 131.935 74.760 132.505 ;
        RECT 74.930 132.395 76.055 132.565 ;
        RECT 74.930 131.765 75.255 132.225 ;
        RECT 75.775 131.935 76.055 132.395 ;
        RECT 76.245 131.935 76.645 132.735 ;
        RECT 76.815 133.465 77.770 133.685 ;
        RECT 78.055 133.645 78.315 134.145 ;
        RECT 78.485 133.815 78.815 134.315 ;
        RECT 78.985 133.725 79.205 134.145 ;
        RECT 79.425 133.815 79.755 134.315 ;
        RECT 78.055 133.475 78.805 133.645 ;
        RECT 76.815 132.565 77.025 133.465 ;
        RECT 77.195 132.735 77.885 133.295 ;
        RECT 78.055 132.655 78.405 133.305 ;
        RECT 76.815 132.395 77.770 132.565 ;
        RECT 78.575 132.485 78.805 133.475 ;
        RECT 77.045 131.765 77.315 132.225 ;
        RECT 77.485 131.935 77.770 132.395 ;
        RECT 78.055 132.315 78.805 132.485 ;
        RECT 78.055 132.025 78.315 132.315 ;
        RECT 78.975 132.245 79.205 133.725 ;
        RECT 79.925 133.645 80.095 134.145 ;
        RECT 80.330 133.930 81.160 134.100 ;
        RECT 81.400 133.935 81.780 134.315 ;
        RECT 79.400 133.475 80.095 133.645 ;
        RECT 79.400 132.505 79.570 133.475 ;
        RECT 79.740 132.685 80.150 133.305 ;
        RECT 80.320 133.255 80.820 133.635 ;
        RECT 79.400 132.315 80.095 132.505 ;
        RECT 80.320 132.385 80.540 133.255 ;
        RECT 80.990 133.085 81.160 133.930 ;
        RECT 81.960 133.765 82.130 134.055 ;
        RECT 82.300 133.935 82.630 134.315 ;
        RECT 83.080 133.845 83.710 134.095 ;
        RECT 83.890 133.935 84.310 134.315 ;
        RECT 83.540 133.765 83.710 133.845 ;
        RECT 84.510 133.765 84.750 134.055 ;
        RECT 81.330 133.515 82.680 133.765 ;
        RECT 81.330 133.255 81.580 133.515 ;
        RECT 82.090 133.085 82.340 133.245 ;
        RECT 80.990 132.915 82.340 133.085 ;
        RECT 80.990 132.875 81.410 132.915 ;
        RECT 80.720 132.325 81.070 132.695 ;
        RECT 78.485 131.765 78.815 132.145 ;
        RECT 78.985 132.025 79.205 132.245 ;
        RECT 79.425 131.765 79.755 132.145 ;
        RECT 79.925 131.985 80.095 132.315 ;
        RECT 81.240 132.145 81.410 132.875 ;
        RECT 82.510 132.745 82.680 133.515 ;
        RECT 81.580 132.415 81.990 132.745 ;
        RECT 82.280 132.405 82.680 132.745 ;
        RECT 82.850 133.335 83.370 133.645 ;
        RECT 83.540 133.595 84.750 133.765 ;
        RECT 84.980 133.625 85.310 134.315 ;
        RECT 82.850 132.575 83.020 133.335 ;
        RECT 83.190 132.745 83.370 133.155 ;
        RECT 83.540 133.085 83.710 133.595 ;
        RECT 85.480 133.445 85.650 134.055 ;
        RECT 85.940 133.595 86.270 134.105 ;
        RECT 85.480 133.425 85.850 133.445 ;
        RECT 83.880 133.255 85.850 133.425 ;
        RECT 83.540 132.915 85.460 133.085 ;
        RECT 83.770 132.575 84.120 132.695 ;
        RECT 82.850 132.405 84.120 132.575 ;
        RECT 80.395 131.945 81.410 132.145 ;
        RECT 81.580 131.765 81.990 132.205 ;
        RECT 82.280 131.975 82.530 132.405 ;
        RECT 82.730 131.765 83.050 132.225 ;
        RECT 84.290 132.155 84.460 132.915 ;
        RECT 85.110 132.855 85.460 132.915 ;
        RECT 84.630 132.685 84.980 132.745 ;
        RECT 84.630 132.415 85.310 132.685 ;
        RECT 85.660 132.360 85.850 133.255 ;
        RECT 83.610 131.985 84.460 132.155 ;
        RECT 84.660 131.765 85.300 132.245 ;
        RECT 85.500 132.030 85.850 132.360 ;
        RECT 86.020 133.005 86.270 133.595 ;
        RECT 86.440 133.175 86.610 134.315 ;
        RECT 86.780 133.295 87.110 134.140 ;
        RECT 87.280 133.465 87.545 134.315 ;
        RECT 86.780 133.175 87.545 133.295 ;
        RECT 87.715 133.225 89.385 134.315 ;
        RECT 86.945 133.125 87.545 133.175 ;
        RECT 86.020 132.675 86.820 133.005 ;
        RECT 86.020 132.025 86.190 132.675 ;
        RECT 86.990 132.575 87.545 133.125 ;
        RECT 86.960 132.535 87.545 132.575 ;
        RECT 86.945 132.505 87.545 132.535 ;
        RECT 86.360 131.765 86.690 132.505 ;
        RECT 86.860 132.445 87.545 132.505 ;
        RECT 87.715 132.535 88.465 133.055 ;
        RECT 88.635 132.705 89.385 133.225 ;
        RECT 89.595 133.175 89.825 134.315 ;
        RECT 89.995 133.165 90.325 134.145 ;
        RECT 90.495 133.175 90.705 134.315 ;
        RECT 90.935 133.880 96.280 134.315 ;
        RECT 89.575 132.755 89.905 133.005 ;
        RECT 86.860 131.945 87.105 132.445 ;
        RECT 87.275 131.765 87.545 132.275 ;
        RECT 87.715 131.765 89.385 132.535 ;
        RECT 89.595 131.765 89.825 132.585 ;
        RECT 90.075 132.565 90.325 133.165 ;
        RECT 89.995 131.935 90.325 132.565 ;
        RECT 90.495 131.765 90.705 132.585 ;
        RECT 92.520 132.310 92.860 133.140 ;
        RECT 94.340 132.630 94.690 133.880 ;
        RECT 96.455 133.225 99.045 134.315 ;
        RECT 96.455 132.535 97.665 133.055 ;
        RECT 97.835 132.705 99.045 133.225 ;
        RECT 99.675 133.150 99.965 134.315 ;
        RECT 100.135 133.880 105.480 134.315 ;
        RECT 90.935 131.765 96.280 132.310 ;
        RECT 96.455 131.765 99.045 132.535 ;
        RECT 99.675 131.765 99.965 132.490 ;
        RECT 101.720 132.310 102.060 133.140 ;
        RECT 103.540 132.630 103.890 133.880 ;
        RECT 105.655 133.225 107.325 134.315 ;
        RECT 105.655 132.535 106.405 133.055 ;
        RECT 106.575 132.705 107.325 133.225 ;
        RECT 107.955 133.225 109.165 134.315 ;
        RECT 107.955 132.685 108.475 133.225 ;
        RECT 100.135 131.765 105.480 132.310 ;
        RECT 105.655 131.765 107.325 132.535 ;
        RECT 108.645 132.515 109.165 133.055 ;
        RECT 107.955 131.765 109.165 132.515 ;
        RECT 35.190 131.595 109.250 131.765 ;
        RECT 35.275 130.845 36.485 131.595 ;
        RECT 36.655 131.050 42.000 131.595 ;
        RECT 42.175 131.050 47.520 131.595 ;
        RECT 47.695 131.050 53.040 131.595 ;
        RECT 53.215 131.050 58.560 131.595 ;
        RECT 35.275 130.305 35.795 130.845 ;
        RECT 35.965 130.135 36.485 130.675 ;
        RECT 38.240 130.220 38.580 131.050 ;
        RECT 35.275 129.045 36.485 130.135 ;
        RECT 40.060 129.480 40.410 130.730 ;
        RECT 43.760 130.220 44.100 131.050 ;
        RECT 45.580 129.480 45.930 130.730 ;
        RECT 49.280 130.220 49.620 131.050 ;
        RECT 51.100 129.480 51.450 130.730 ;
        RECT 54.800 130.220 55.140 131.050 ;
        RECT 58.735 130.825 60.405 131.595 ;
        RECT 61.035 130.870 61.325 131.595 ;
        RECT 61.495 130.825 63.165 131.595 ;
        RECT 63.795 130.855 64.180 131.425 ;
        RECT 64.350 131.135 64.675 131.595 ;
        RECT 65.195 130.965 65.475 131.425 ;
        RECT 56.620 129.480 56.970 130.730 ;
        RECT 58.735 130.305 59.485 130.825 ;
        RECT 59.655 130.135 60.405 130.655 ;
        RECT 61.495 130.305 62.245 130.825 ;
        RECT 36.655 129.045 42.000 129.480 ;
        RECT 42.175 129.045 47.520 129.480 ;
        RECT 47.695 129.045 53.040 129.480 ;
        RECT 53.215 129.045 58.560 129.480 ;
        RECT 58.735 129.045 60.405 130.135 ;
        RECT 61.035 129.045 61.325 130.210 ;
        RECT 62.415 130.135 63.165 130.655 ;
        RECT 61.495 129.045 63.165 130.135 ;
        RECT 63.795 130.185 64.075 130.855 ;
        RECT 64.350 130.795 65.475 130.965 ;
        RECT 64.350 130.685 64.800 130.795 ;
        RECT 64.245 130.355 64.800 130.685 ;
        RECT 65.665 130.625 66.065 131.425 ;
        RECT 66.465 131.135 66.735 131.595 ;
        RECT 66.905 130.965 67.190 131.425 ;
        RECT 63.795 129.215 64.180 130.185 ;
        RECT 64.350 129.895 64.800 130.355 ;
        RECT 64.970 130.065 66.065 130.625 ;
        RECT 64.350 129.675 65.475 129.895 ;
        RECT 64.350 129.045 64.675 129.505 ;
        RECT 65.195 129.215 65.475 129.675 ;
        RECT 65.665 129.215 66.065 130.065 ;
        RECT 66.235 130.795 67.190 130.965 ;
        RECT 67.475 130.845 68.685 131.595 ;
        RECT 68.855 131.085 69.125 131.595 ;
        RECT 69.295 130.915 69.540 131.415 ;
        RECT 68.855 130.855 69.540 130.915 ;
        RECT 69.710 130.855 70.040 131.595 ;
        RECT 66.235 129.895 66.445 130.795 ;
        RECT 66.615 130.065 67.305 130.625 ;
        RECT 67.475 130.305 67.995 130.845 ;
        RECT 68.855 130.825 69.455 130.855 ;
        RECT 68.855 130.785 69.440 130.825 ;
        RECT 68.165 130.135 68.685 130.675 ;
        RECT 66.235 129.675 67.190 129.895 ;
        RECT 66.465 129.045 66.735 129.505 ;
        RECT 66.905 129.215 67.190 129.675 ;
        RECT 67.475 129.045 68.685 130.135 ;
        RECT 68.855 130.235 69.410 130.785 ;
        RECT 70.210 130.685 70.380 131.335 ;
        RECT 69.580 130.355 70.380 130.685 ;
        RECT 68.855 130.185 69.455 130.235 ;
        RECT 68.855 130.065 69.620 130.185 ;
        RECT 68.855 129.045 69.120 129.895 ;
        RECT 69.290 129.220 69.620 130.065 ;
        RECT 69.790 129.045 69.960 130.185 ;
        RECT 70.130 129.765 70.380 130.355 ;
        RECT 70.550 131.000 70.900 131.330 ;
        RECT 71.100 131.115 71.740 131.595 ;
        RECT 71.940 131.205 72.790 131.375 ;
        RECT 70.550 130.105 70.740 131.000 ;
        RECT 71.090 130.675 71.770 130.945 ;
        RECT 71.420 130.615 71.770 130.675 ;
        RECT 70.940 130.445 71.290 130.505 ;
        RECT 71.940 130.445 72.110 131.205 ;
        RECT 73.350 131.135 73.670 131.595 ;
        RECT 73.870 130.955 74.120 131.385 ;
        RECT 74.410 131.155 74.820 131.595 ;
        RECT 74.990 131.215 76.005 131.415 ;
        RECT 72.280 130.785 73.550 130.955 ;
        RECT 72.280 130.665 72.630 130.785 ;
        RECT 70.940 130.275 72.860 130.445 ;
        RECT 70.550 129.935 72.520 130.105 ;
        RECT 70.550 129.915 70.920 129.935 ;
        RECT 70.130 129.255 70.460 129.765 ;
        RECT 70.750 129.305 70.920 129.915 ;
        RECT 72.690 129.765 72.860 130.275 ;
        RECT 73.030 130.205 73.210 130.615 ;
        RECT 73.380 130.025 73.550 130.785 ;
        RECT 71.090 129.045 71.420 129.735 ;
        RECT 71.650 129.595 72.860 129.765 ;
        RECT 73.030 129.715 73.550 130.025 ;
        RECT 73.720 130.615 74.120 130.955 ;
        RECT 74.410 130.615 74.820 130.945 ;
        RECT 73.720 129.845 73.890 130.615 ;
        RECT 74.990 130.485 75.160 131.215 ;
        RECT 76.305 131.045 76.475 131.375 ;
        RECT 76.645 131.215 76.975 131.595 ;
        RECT 77.195 131.115 77.415 131.335 ;
        RECT 77.585 131.215 77.915 131.595 ;
        RECT 75.330 130.665 75.680 131.035 ;
        RECT 74.990 130.445 75.410 130.485 ;
        RECT 74.060 130.275 75.410 130.445 ;
        RECT 74.060 130.115 74.310 130.275 ;
        RECT 74.820 129.845 75.070 130.105 ;
        RECT 73.720 129.595 75.070 129.845 ;
        RECT 71.650 129.305 71.890 129.595 ;
        RECT 72.690 129.515 72.860 129.595 ;
        RECT 72.090 129.045 72.510 129.425 ;
        RECT 72.690 129.265 73.320 129.515 ;
        RECT 73.770 129.045 74.100 129.425 ;
        RECT 74.270 129.305 74.440 129.595 ;
        RECT 75.240 129.430 75.410 130.275 ;
        RECT 75.860 130.105 76.080 130.975 ;
        RECT 76.305 130.855 77.000 131.045 ;
        RECT 75.580 129.725 76.080 130.105 ;
        RECT 76.250 130.055 76.660 130.675 ;
        RECT 76.830 129.885 77.000 130.855 ;
        RECT 76.305 129.715 77.000 129.885 ;
        RECT 74.620 129.045 75.000 129.425 ;
        RECT 75.240 129.260 76.070 129.430 ;
        RECT 76.305 129.215 76.475 129.715 ;
        RECT 77.195 129.635 77.425 131.115 ;
        RECT 78.085 131.045 78.345 131.335 ;
        RECT 77.595 130.875 78.345 131.045 ;
        RECT 77.595 129.885 77.825 130.875 ;
        RECT 78.515 130.825 82.025 131.595 ;
        RECT 77.995 130.055 78.345 130.705 ;
        RECT 78.515 130.305 80.165 130.825 ;
        RECT 83.175 130.775 83.385 131.595 ;
        RECT 83.555 130.795 83.885 131.425 ;
        RECT 80.335 130.135 82.025 130.655 ;
        RECT 83.555 130.195 83.805 130.795 ;
        RECT 84.055 130.775 84.285 131.595 ;
        RECT 84.495 130.825 86.165 131.595 ;
        RECT 86.795 130.870 87.085 131.595 ;
        RECT 87.255 131.050 92.600 131.595 ;
        RECT 92.775 131.050 98.120 131.595 ;
        RECT 98.295 131.050 103.640 131.595 ;
        RECT 83.975 130.355 84.305 130.605 ;
        RECT 84.495 130.305 85.245 130.825 ;
        RECT 77.595 129.715 78.345 129.885 ;
        RECT 76.645 129.045 76.975 129.545 ;
        RECT 77.195 129.215 77.415 129.635 ;
        RECT 77.585 129.045 77.915 129.545 ;
        RECT 78.085 129.215 78.345 129.715 ;
        RECT 78.515 129.045 82.025 130.135 ;
        RECT 83.175 129.045 83.385 130.185 ;
        RECT 83.555 129.215 83.885 130.195 ;
        RECT 84.055 129.045 84.285 130.185 ;
        RECT 85.415 130.135 86.165 130.655 ;
        RECT 88.840 130.220 89.180 131.050 ;
        RECT 84.495 129.045 86.165 130.135 ;
        RECT 86.795 129.045 87.085 130.210 ;
        RECT 90.660 129.480 91.010 130.730 ;
        RECT 94.360 130.220 94.700 131.050 ;
        RECT 96.180 129.480 96.530 130.730 ;
        RECT 99.880 130.220 100.220 131.050 ;
        RECT 103.815 130.825 107.325 131.595 ;
        RECT 107.955 130.845 109.165 131.595 ;
        RECT 101.700 129.480 102.050 130.730 ;
        RECT 103.815 130.305 105.465 130.825 ;
        RECT 105.635 130.135 107.325 130.655 ;
        RECT 87.255 129.045 92.600 129.480 ;
        RECT 92.775 129.045 98.120 129.480 ;
        RECT 98.295 129.045 103.640 129.480 ;
        RECT 103.815 129.045 107.325 130.135 ;
        RECT 107.955 130.135 108.475 130.675 ;
        RECT 108.645 130.305 109.165 130.845 ;
        RECT 107.955 129.045 109.165 130.135 ;
        RECT 35.190 128.875 109.250 129.045 ;
        RECT 35.275 127.785 36.485 128.875 ;
        RECT 36.655 128.440 42.000 128.875 ;
        RECT 42.175 128.440 47.520 128.875 ;
        RECT 35.275 127.075 35.795 127.615 ;
        RECT 35.965 127.245 36.485 127.785 ;
        RECT 35.275 126.325 36.485 127.075 ;
        RECT 38.240 126.870 38.580 127.700 ;
        RECT 40.060 127.190 40.410 128.440 ;
        RECT 43.760 126.870 44.100 127.700 ;
        RECT 45.580 127.190 45.930 128.440 ;
        RECT 48.155 127.710 48.445 128.875 ;
        RECT 48.615 128.440 53.960 128.875 ;
        RECT 54.135 128.440 59.480 128.875 ;
        RECT 36.655 126.325 42.000 126.870 ;
        RECT 42.175 126.325 47.520 126.870 ;
        RECT 48.155 126.325 48.445 127.050 ;
        RECT 50.200 126.870 50.540 127.700 ;
        RECT 52.020 127.190 52.370 128.440 ;
        RECT 55.720 126.870 56.060 127.700 ;
        RECT 57.540 127.190 57.890 128.440 ;
        RECT 59.655 127.785 63.165 128.875 ;
        RECT 59.655 127.095 61.305 127.615 ;
        RECT 61.475 127.265 63.165 127.785 ;
        RECT 63.795 127.270 64.075 128.705 ;
        RECT 64.245 128.100 64.955 128.875 ;
        RECT 65.125 127.930 65.455 128.705 ;
        RECT 64.305 127.715 65.455 127.930 ;
        RECT 48.615 126.325 53.960 126.870 ;
        RECT 54.135 126.325 59.480 126.870 ;
        RECT 59.655 126.325 63.165 127.095 ;
        RECT 63.795 126.495 64.135 127.270 ;
        RECT 64.305 127.145 64.590 127.715 ;
        RECT 64.775 127.315 65.245 127.545 ;
        RECT 65.650 127.515 65.865 128.630 ;
        RECT 66.045 128.155 66.375 128.875 ;
        RECT 66.555 128.440 71.900 128.875 ;
        RECT 66.155 127.515 66.385 127.855 ;
        RECT 65.415 127.335 65.865 127.515 ;
        RECT 65.415 127.315 65.745 127.335 ;
        RECT 66.055 127.315 66.385 127.515 ;
        RECT 64.305 126.955 65.015 127.145 ;
        RECT 64.715 126.815 65.015 126.955 ;
        RECT 65.205 126.955 66.385 127.145 ;
        RECT 65.205 126.875 65.535 126.955 ;
        RECT 64.715 126.805 65.030 126.815 ;
        RECT 64.715 126.795 65.040 126.805 ;
        RECT 64.715 126.790 65.050 126.795 ;
        RECT 64.305 126.325 64.475 126.785 ;
        RECT 64.715 126.780 65.055 126.790 ;
        RECT 64.715 126.775 65.060 126.780 ;
        RECT 64.715 126.765 65.065 126.775 ;
        RECT 64.715 126.760 65.070 126.765 ;
        RECT 64.715 126.495 65.075 126.760 ;
        RECT 65.705 126.325 65.875 126.785 ;
        RECT 66.045 126.495 66.385 126.955 ;
        RECT 68.140 126.870 68.480 127.700 ;
        RECT 69.960 127.190 70.310 128.440 ;
        RECT 72.075 127.785 73.745 128.875 ;
        RECT 72.075 127.095 72.825 127.615 ;
        RECT 72.995 127.265 73.745 127.785 ;
        RECT 73.915 127.710 74.205 128.875 ;
        RECT 74.375 128.440 79.720 128.875 ;
        RECT 79.895 128.440 85.240 128.875 ;
        RECT 85.415 128.440 90.760 128.875 ;
        RECT 90.935 128.440 96.280 128.875 ;
        RECT 66.555 126.325 71.900 126.870 ;
        RECT 72.075 126.325 73.745 127.095 ;
        RECT 73.915 126.325 74.205 127.050 ;
        RECT 75.960 126.870 76.300 127.700 ;
        RECT 77.780 127.190 78.130 128.440 ;
        RECT 81.480 126.870 81.820 127.700 ;
        RECT 83.300 127.190 83.650 128.440 ;
        RECT 87.000 126.870 87.340 127.700 ;
        RECT 88.820 127.190 89.170 128.440 ;
        RECT 92.520 126.870 92.860 127.700 ;
        RECT 94.340 127.190 94.690 128.440 ;
        RECT 96.455 127.785 99.045 128.875 ;
        RECT 96.455 127.095 97.665 127.615 ;
        RECT 97.835 127.265 99.045 127.785 ;
        RECT 99.675 127.710 99.965 128.875 ;
        RECT 100.135 128.440 105.480 128.875 ;
        RECT 74.375 126.325 79.720 126.870 ;
        RECT 79.895 126.325 85.240 126.870 ;
        RECT 85.415 126.325 90.760 126.870 ;
        RECT 90.935 126.325 96.280 126.870 ;
        RECT 96.455 126.325 99.045 127.095 ;
        RECT 99.675 126.325 99.965 127.050 ;
        RECT 101.720 126.870 102.060 127.700 ;
        RECT 103.540 127.190 103.890 128.440 ;
        RECT 105.655 127.785 107.325 128.875 ;
        RECT 105.655 127.095 106.405 127.615 ;
        RECT 106.575 127.265 107.325 127.785 ;
        RECT 107.955 127.785 109.165 128.875 ;
        RECT 107.955 127.245 108.475 127.785 ;
        RECT 100.135 126.325 105.480 126.870 ;
        RECT 105.655 126.325 107.325 127.095 ;
        RECT 108.645 127.075 109.165 127.615 ;
        RECT 107.955 126.325 109.165 127.075 ;
        RECT 35.190 126.155 109.250 126.325 ;
        RECT 35.275 125.405 36.485 126.155 ;
        RECT 36.655 125.610 42.000 126.155 ;
        RECT 42.175 125.610 47.520 126.155 ;
        RECT 47.695 125.610 53.040 126.155 ;
        RECT 53.215 125.610 58.560 126.155 ;
        RECT 35.275 124.865 35.795 125.405 ;
        RECT 35.965 124.695 36.485 125.235 ;
        RECT 38.240 124.780 38.580 125.610 ;
        RECT 35.275 123.605 36.485 124.695 ;
        RECT 40.060 124.040 40.410 125.290 ;
        RECT 43.760 124.780 44.100 125.610 ;
        RECT 45.580 124.040 45.930 125.290 ;
        RECT 49.280 124.780 49.620 125.610 ;
        RECT 51.100 124.040 51.450 125.290 ;
        RECT 54.800 124.780 55.140 125.610 ;
        RECT 58.735 125.385 60.405 126.155 ;
        RECT 61.035 125.430 61.325 126.155 ;
        RECT 61.495 125.610 66.840 126.155 ;
        RECT 67.015 125.610 72.360 126.155 ;
        RECT 72.535 125.610 77.880 126.155 ;
        RECT 78.055 125.610 83.400 126.155 ;
        RECT 56.620 124.040 56.970 125.290 ;
        RECT 58.735 124.865 59.485 125.385 ;
        RECT 59.655 124.695 60.405 125.215 ;
        RECT 63.080 124.780 63.420 125.610 ;
        RECT 36.655 123.605 42.000 124.040 ;
        RECT 42.175 123.605 47.520 124.040 ;
        RECT 47.695 123.605 53.040 124.040 ;
        RECT 53.215 123.605 58.560 124.040 ;
        RECT 58.735 123.605 60.405 124.695 ;
        RECT 61.035 123.605 61.325 124.770 ;
        RECT 64.900 124.040 65.250 125.290 ;
        RECT 68.600 124.780 68.940 125.610 ;
        RECT 70.420 124.040 70.770 125.290 ;
        RECT 74.120 124.780 74.460 125.610 ;
        RECT 75.940 124.040 76.290 125.290 ;
        RECT 79.640 124.780 79.980 125.610 ;
        RECT 83.575 125.385 86.165 126.155 ;
        RECT 86.795 125.430 87.085 126.155 ;
        RECT 87.255 125.610 92.600 126.155 ;
        RECT 92.775 125.610 98.120 126.155 ;
        RECT 98.295 125.610 103.640 126.155 ;
        RECT 81.460 124.040 81.810 125.290 ;
        RECT 83.575 124.865 84.785 125.385 ;
        RECT 84.955 124.695 86.165 125.215 ;
        RECT 88.840 124.780 89.180 125.610 ;
        RECT 61.495 123.605 66.840 124.040 ;
        RECT 67.015 123.605 72.360 124.040 ;
        RECT 72.535 123.605 77.880 124.040 ;
        RECT 78.055 123.605 83.400 124.040 ;
        RECT 83.575 123.605 86.165 124.695 ;
        RECT 86.795 123.605 87.085 124.770 ;
        RECT 90.660 124.040 91.010 125.290 ;
        RECT 94.360 124.780 94.700 125.610 ;
        RECT 96.180 124.040 96.530 125.290 ;
        RECT 99.880 124.780 100.220 125.610 ;
        RECT 103.815 125.385 107.325 126.155 ;
        RECT 107.955 125.405 109.165 126.155 ;
        RECT 101.700 124.040 102.050 125.290 ;
        RECT 103.815 124.865 105.465 125.385 ;
        RECT 105.635 124.695 107.325 125.215 ;
        RECT 87.255 123.605 92.600 124.040 ;
        RECT 92.775 123.605 98.120 124.040 ;
        RECT 98.295 123.605 103.640 124.040 ;
        RECT 103.815 123.605 107.325 124.695 ;
        RECT 107.955 124.695 108.475 125.235 ;
        RECT 108.645 124.865 109.165 125.405 ;
        RECT 107.955 123.605 109.165 124.695 ;
        RECT 35.190 123.435 109.250 123.605 ;
        RECT 35.275 122.345 36.485 123.435 ;
        RECT 36.655 123.000 42.000 123.435 ;
        RECT 42.175 123.000 47.520 123.435 ;
        RECT 35.275 121.635 35.795 122.175 ;
        RECT 35.965 121.805 36.485 122.345 ;
        RECT 35.275 120.885 36.485 121.635 ;
        RECT 38.240 121.430 38.580 122.260 ;
        RECT 40.060 121.750 40.410 123.000 ;
        RECT 43.760 121.430 44.100 122.260 ;
        RECT 45.580 121.750 45.930 123.000 ;
        RECT 48.155 122.270 48.445 123.435 ;
        RECT 48.615 123.000 53.960 123.435 ;
        RECT 54.135 123.000 59.480 123.435 ;
        RECT 59.655 123.000 65.000 123.435 ;
        RECT 65.175 123.000 70.520 123.435 ;
        RECT 36.655 120.885 42.000 121.430 ;
        RECT 42.175 120.885 47.520 121.430 ;
        RECT 48.155 120.885 48.445 121.610 ;
        RECT 50.200 121.430 50.540 122.260 ;
        RECT 52.020 121.750 52.370 123.000 ;
        RECT 55.720 121.430 56.060 122.260 ;
        RECT 57.540 121.750 57.890 123.000 ;
        RECT 61.240 121.430 61.580 122.260 ;
        RECT 63.060 121.750 63.410 123.000 ;
        RECT 66.760 121.430 67.100 122.260 ;
        RECT 68.580 121.750 68.930 123.000 ;
        RECT 70.695 122.345 73.285 123.435 ;
        RECT 70.695 121.655 71.905 122.175 ;
        RECT 72.075 121.825 73.285 122.345 ;
        RECT 73.915 122.270 74.205 123.435 ;
        RECT 74.375 123.000 79.720 123.435 ;
        RECT 79.895 123.000 85.240 123.435 ;
        RECT 85.415 123.000 90.760 123.435 ;
        RECT 90.935 123.000 96.280 123.435 ;
        RECT 48.615 120.885 53.960 121.430 ;
        RECT 54.135 120.885 59.480 121.430 ;
        RECT 59.655 120.885 65.000 121.430 ;
        RECT 65.175 120.885 70.520 121.430 ;
        RECT 70.695 120.885 73.285 121.655 ;
        RECT 73.915 120.885 74.205 121.610 ;
        RECT 75.960 121.430 76.300 122.260 ;
        RECT 77.780 121.750 78.130 123.000 ;
        RECT 81.480 121.430 81.820 122.260 ;
        RECT 83.300 121.750 83.650 123.000 ;
        RECT 87.000 121.430 87.340 122.260 ;
        RECT 88.820 121.750 89.170 123.000 ;
        RECT 92.520 121.430 92.860 122.260 ;
        RECT 94.340 121.750 94.690 123.000 ;
        RECT 96.455 122.345 99.045 123.435 ;
        RECT 96.455 121.655 97.665 122.175 ;
        RECT 97.835 121.825 99.045 122.345 ;
        RECT 99.675 122.270 99.965 123.435 ;
        RECT 100.135 123.000 105.480 123.435 ;
        RECT 74.375 120.885 79.720 121.430 ;
        RECT 79.895 120.885 85.240 121.430 ;
        RECT 85.415 120.885 90.760 121.430 ;
        RECT 90.935 120.885 96.280 121.430 ;
        RECT 96.455 120.885 99.045 121.655 ;
        RECT 99.675 120.885 99.965 121.610 ;
        RECT 101.720 121.430 102.060 122.260 ;
        RECT 103.540 121.750 103.890 123.000 ;
        RECT 105.655 122.345 107.325 123.435 ;
        RECT 105.655 121.655 106.405 122.175 ;
        RECT 106.575 121.825 107.325 122.345 ;
        RECT 107.955 122.345 109.165 123.435 ;
        RECT 107.955 121.805 108.475 122.345 ;
        RECT 100.135 120.885 105.480 121.430 ;
        RECT 105.655 120.885 107.325 121.655 ;
        RECT 108.645 121.635 109.165 122.175 ;
        RECT 107.955 120.885 109.165 121.635 ;
        RECT 35.190 120.715 109.250 120.885 ;
        RECT 35.275 119.965 36.485 120.715 ;
        RECT 36.655 120.170 42.000 120.715 ;
        RECT 42.175 120.170 47.520 120.715 ;
        RECT 47.695 120.170 53.040 120.715 ;
        RECT 53.215 120.170 58.560 120.715 ;
        RECT 35.275 119.425 35.795 119.965 ;
        RECT 35.965 119.255 36.485 119.795 ;
        RECT 38.240 119.340 38.580 120.170 ;
        RECT 35.275 118.165 36.485 119.255 ;
        RECT 40.060 118.600 40.410 119.850 ;
        RECT 43.760 119.340 44.100 120.170 ;
        RECT 45.580 118.600 45.930 119.850 ;
        RECT 49.280 119.340 49.620 120.170 ;
        RECT 51.100 118.600 51.450 119.850 ;
        RECT 54.800 119.340 55.140 120.170 ;
        RECT 58.735 119.945 60.405 120.715 ;
        RECT 61.035 119.990 61.325 120.715 ;
        RECT 61.495 120.170 66.840 120.715 ;
        RECT 67.015 120.170 72.360 120.715 ;
        RECT 72.535 120.170 77.880 120.715 ;
        RECT 78.055 120.170 83.400 120.715 ;
        RECT 56.620 118.600 56.970 119.850 ;
        RECT 58.735 119.425 59.485 119.945 ;
        RECT 59.655 119.255 60.405 119.775 ;
        RECT 63.080 119.340 63.420 120.170 ;
        RECT 36.655 118.165 42.000 118.600 ;
        RECT 42.175 118.165 47.520 118.600 ;
        RECT 47.695 118.165 53.040 118.600 ;
        RECT 53.215 118.165 58.560 118.600 ;
        RECT 58.735 118.165 60.405 119.255 ;
        RECT 61.035 118.165 61.325 119.330 ;
        RECT 64.900 118.600 65.250 119.850 ;
        RECT 68.600 119.340 68.940 120.170 ;
        RECT 70.420 118.600 70.770 119.850 ;
        RECT 74.120 119.340 74.460 120.170 ;
        RECT 75.940 118.600 76.290 119.850 ;
        RECT 79.640 119.340 79.980 120.170 ;
        RECT 83.575 119.945 86.165 120.715 ;
        RECT 86.795 119.990 87.085 120.715 ;
        RECT 87.255 120.170 92.600 120.715 ;
        RECT 92.775 120.170 98.120 120.715 ;
        RECT 98.295 120.170 103.640 120.715 ;
        RECT 81.460 118.600 81.810 119.850 ;
        RECT 83.575 119.425 84.785 119.945 ;
        RECT 84.955 119.255 86.165 119.775 ;
        RECT 88.840 119.340 89.180 120.170 ;
        RECT 61.495 118.165 66.840 118.600 ;
        RECT 67.015 118.165 72.360 118.600 ;
        RECT 72.535 118.165 77.880 118.600 ;
        RECT 78.055 118.165 83.400 118.600 ;
        RECT 83.575 118.165 86.165 119.255 ;
        RECT 86.795 118.165 87.085 119.330 ;
        RECT 90.660 118.600 91.010 119.850 ;
        RECT 94.360 119.340 94.700 120.170 ;
        RECT 96.180 118.600 96.530 119.850 ;
        RECT 99.880 119.340 100.220 120.170 ;
        RECT 103.815 119.945 107.325 120.715 ;
        RECT 107.955 119.965 109.165 120.715 ;
        RECT 101.700 118.600 102.050 119.850 ;
        RECT 103.815 119.425 105.465 119.945 ;
        RECT 105.635 119.255 107.325 119.775 ;
        RECT 87.255 118.165 92.600 118.600 ;
        RECT 92.775 118.165 98.120 118.600 ;
        RECT 98.295 118.165 103.640 118.600 ;
        RECT 103.815 118.165 107.325 119.255 ;
        RECT 107.955 119.255 108.475 119.795 ;
        RECT 108.645 119.425 109.165 119.965 ;
        RECT 107.955 118.165 109.165 119.255 ;
        RECT 35.190 117.995 109.250 118.165 ;
        RECT 35.275 116.905 36.485 117.995 ;
        RECT 36.655 117.560 42.000 117.995 ;
        RECT 42.175 117.560 47.520 117.995 ;
        RECT 35.275 116.195 35.795 116.735 ;
        RECT 35.965 116.365 36.485 116.905 ;
        RECT 35.275 115.445 36.485 116.195 ;
        RECT 38.240 115.990 38.580 116.820 ;
        RECT 40.060 116.310 40.410 117.560 ;
        RECT 43.760 115.990 44.100 116.820 ;
        RECT 45.580 116.310 45.930 117.560 ;
        RECT 48.155 116.830 48.445 117.995 ;
        RECT 48.615 117.560 53.960 117.995 ;
        RECT 54.135 117.560 59.480 117.995 ;
        RECT 59.655 117.560 65.000 117.995 ;
        RECT 65.175 117.560 70.520 117.995 ;
        RECT 36.655 115.445 42.000 115.990 ;
        RECT 42.175 115.445 47.520 115.990 ;
        RECT 48.155 115.445 48.445 116.170 ;
        RECT 50.200 115.990 50.540 116.820 ;
        RECT 52.020 116.310 52.370 117.560 ;
        RECT 55.720 115.990 56.060 116.820 ;
        RECT 57.540 116.310 57.890 117.560 ;
        RECT 61.240 115.990 61.580 116.820 ;
        RECT 63.060 116.310 63.410 117.560 ;
        RECT 66.760 115.990 67.100 116.820 ;
        RECT 68.580 116.310 68.930 117.560 ;
        RECT 70.695 116.905 73.285 117.995 ;
        RECT 70.695 116.215 71.905 116.735 ;
        RECT 72.075 116.385 73.285 116.905 ;
        RECT 73.915 116.830 74.205 117.995 ;
        RECT 74.375 117.560 79.720 117.995 ;
        RECT 79.895 117.560 85.240 117.995 ;
        RECT 85.415 117.560 90.760 117.995 ;
        RECT 90.935 117.560 96.280 117.995 ;
        RECT 48.615 115.445 53.960 115.990 ;
        RECT 54.135 115.445 59.480 115.990 ;
        RECT 59.655 115.445 65.000 115.990 ;
        RECT 65.175 115.445 70.520 115.990 ;
        RECT 70.695 115.445 73.285 116.215 ;
        RECT 73.915 115.445 74.205 116.170 ;
        RECT 75.960 115.990 76.300 116.820 ;
        RECT 77.780 116.310 78.130 117.560 ;
        RECT 81.480 115.990 81.820 116.820 ;
        RECT 83.300 116.310 83.650 117.560 ;
        RECT 87.000 115.990 87.340 116.820 ;
        RECT 88.820 116.310 89.170 117.560 ;
        RECT 92.520 115.990 92.860 116.820 ;
        RECT 94.340 116.310 94.690 117.560 ;
        RECT 96.455 116.905 99.045 117.995 ;
        RECT 96.455 116.215 97.665 116.735 ;
        RECT 97.835 116.385 99.045 116.905 ;
        RECT 99.675 116.830 99.965 117.995 ;
        RECT 100.135 117.560 105.480 117.995 ;
        RECT 74.375 115.445 79.720 115.990 ;
        RECT 79.895 115.445 85.240 115.990 ;
        RECT 85.415 115.445 90.760 115.990 ;
        RECT 90.935 115.445 96.280 115.990 ;
        RECT 96.455 115.445 99.045 116.215 ;
        RECT 99.675 115.445 99.965 116.170 ;
        RECT 101.720 115.990 102.060 116.820 ;
        RECT 103.540 116.310 103.890 117.560 ;
        RECT 105.655 116.905 107.325 117.995 ;
        RECT 105.655 116.215 106.405 116.735 ;
        RECT 106.575 116.385 107.325 116.905 ;
        RECT 107.955 116.905 109.165 117.995 ;
        RECT 107.955 116.365 108.475 116.905 ;
        RECT 100.135 115.445 105.480 115.990 ;
        RECT 105.655 115.445 107.325 116.215 ;
        RECT 108.645 116.195 109.165 116.735 ;
        RECT 107.955 115.445 109.165 116.195 ;
        RECT 35.190 115.275 109.250 115.445 ;
        RECT 35.275 114.525 36.485 115.275 ;
        RECT 36.655 114.730 42.000 115.275 ;
        RECT 42.175 114.730 47.520 115.275 ;
        RECT 47.695 114.730 53.040 115.275 ;
        RECT 53.215 114.730 58.560 115.275 ;
        RECT 35.275 113.985 35.795 114.525 ;
        RECT 35.965 113.815 36.485 114.355 ;
        RECT 38.240 113.900 38.580 114.730 ;
        RECT 35.275 112.725 36.485 113.815 ;
        RECT 40.060 113.160 40.410 114.410 ;
        RECT 43.760 113.900 44.100 114.730 ;
        RECT 45.580 113.160 45.930 114.410 ;
        RECT 49.280 113.900 49.620 114.730 ;
        RECT 51.100 113.160 51.450 114.410 ;
        RECT 54.800 113.900 55.140 114.730 ;
        RECT 58.735 114.505 60.405 115.275 ;
        RECT 61.035 114.550 61.325 115.275 ;
        RECT 61.495 114.730 66.840 115.275 ;
        RECT 67.015 114.730 72.360 115.275 ;
        RECT 72.535 114.730 77.880 115.275 ;
        RECT 78.055 114.730 83.400 115.275 ;
        RECT 56.620 113.160 56.970 114.410 ;
        RECT 58.735 113.985 59.485 114.505 ;
        RECT 59.655 113.815 60.405 114.335 ;
        RECT 63.080 113.900 63.420 114.730 ;
        RECT 36.655 112.725 42.000 113.160 ;
        RECT 42.175 112.725 47.520 113.160 ;
        RECT 47.695 112.725 53.040 113.160 ;
        RECT 53.215 112.725 58.560 113.160 ;
        RECT 58.735 112.725 60.405 113.815 ;
        RECT 61.035 112.725 61.325 113.890 ;
        RECT 64.900 113.160 65.250 114.410 ;
        RECT 68.600 113.900 68.940 114.730 ;
        RECT 70.420 113.160 70.770 114.410 ;
        RECT 74.120 113.900 74.460 114.730 ;
        RECT 75.940 113.160 76.290 114.410 ;
        RECT 79.640 113.900 79.980 114.730 ;
        RECT 83.575 114.505 86.165 115.275 ;
        RECT 86.795 114.550 87.085 115.275 ;
        RECT 87.255 114.730 92.600 115.275 ;
        RECT 92.775 114.730 98.120 115.275 ;
        RECT 98.295 114.730 103.640 115.275 ;
        RECT 81.460 113.160 81.810 114.410 ;
        RECT 83.575 113.985 84.785 114.505 ;
        RECT 84.955 113.815 86.165 114.335 ;
        RECT 88.840 113.900 89.180 114.730 ;
        RECT 61.495 112.725 66.840 113.160 ;
        RECT 67.015 112.725 72.360 113.160 ;
        RECT 72.535 112.725 77.880 113.160 ;
        RECT 78.055 112.725 83.400 113.160 ;
        RECT 83.575 112.725 86.165 113.815 ;
        RECT 86.795 112.725 87.085 113.890 ;
        RECT 90.660 113.160 91.010 114.410 ;
        RECT 94.360 113.900 94.700 114.730 ;
        RECT 96.180 113.160 96.530 114.410 ;
        RECT 99.880 113.900 100.220 114.730 ;
        RECT 103.815 114.505 107.325 115.275 ;
        RECT 107.955 114.525 109.165 115.275 ;
        RECT 101.700 113.160 102.050 114.410 ;
        RECT 103.815 113.985 105.465 114.505 ;
        RECT 105.635 113.815 107.325 114.335 ;
        RECT 87.255 112.725 92.600 113.160 ;
        RECT 92.775 112.725 98.120 113.160 ;
        RECT 98.295 112.725 103.640 113.160 ;
        RECT 103.815 112.725 107.325 113.815 ;
        RECT 107.955 113.815 108.475 114.355 ;
        RECT 108.645 113.985 109.165 114.525 ;
        RECT 107.955 112.725 109.165 113.815 ;
        RECT 35.190 112.555 109.250 112.725 ;
        RECT 35.275 111.465 36.485 112.555 ;
        RECT 36.655 112.120 42.000 112.555 ;
        RECT 42.175 112.120 47.520 112.555 ;
        RECT 35.275 110.755 35.795 111.295 ;
        RECT 35.965 110.925 36.485 111.465 ;
        RECT 35.275 110.005 36.485 110.755 ;
        RECT 38.240 110.550 38.580 111.380 ;
        RECT 40.060 110.870 40.410 112.120 ;
        RECT 43.760 110.550 44.100 111.380 ;
        RECT 45.580 110.870 45.930 112.120 ;
        RECT 48.155 111.390 48.445 112.555 ;
        RECT 48.615 112.120 53.960 112.555 ;
        RECT 54.135 112.120 59.480 112.555 ;
        RECT 59.655 112.120 65.000 112.555 ;
        RECT 65.175 112.120 70.520 112.555 ;
        RECT 36.655 110.005 42.000 110.550 ;
        RECT 42.175 110.005 47.520 110.550 ;
        RECT 48.155 110.005 48.445 110.730 ;
        RECT 50.200 110.550 50.540 111.380 ;
        RECT 52.020 110.870 52.370 112.120 ;
        RECT 55.720 110.550 56.060 111.380 ;
        RECT 57.540 110.870 57.890 112.120 ;
        RECT 61.240 110.550 61.580 111.380 ;
        RECT 63.060 110.870 63.410 112.120 ;
        RECT 66.760 110.550 67.100 111.380 ;
        RECT 68.580 110.870 68.930 112.120 ;
        RECT 70.695 111.465 73.285 112.555 ;
        RECT 70.695 110.775 71.905 111.295 ;
        RECT 72.075 110.945 73.285 111.465 ;
        RECT 73.915 111.390 74.205 112.555 ;
        RECT 74.375 112.120 79.720 112.555 ;
        RECT 79.895 112.120 85.240 112.555 ;
        RECT 85.415 112.120 90.760 112.555 ;
        RECT 90.935 112.120 96.280 112.555 ;
        RECT 48.615 110.005 53.960 110.550 ;
        RECT 54.135 110.005 59.480 110.550 ;
        RECT 59.655 110.005 65.000 110.550 ;
        RECT 65.175 110.005 70.520 110.550 ;
        RECT 70.695 110.005 73.285 110.775 ;
        RECT 73.915 110.005 74.205 110.730 ;
        RECT 75.960 110.550 76.300 111.380 ;
        RECT 77.780 110.870 78.130 112.120 ;
        RECT 81.480 110.550 81.820 111.380 ;
        RECT 83.300 110.870 83.650 112.120 ;
        RECT 87.000 110.550 87.340 111.380 ;
        RECT 88.820 110.870 89.170 112.120 ;
        RECT 92.520 110.550 92.860 111.380 ;
        RECT 94.340 110.870 94.690 112.120 ;
        RECT 96.455 111.465 99.045 112.555 ;
        RECT 96.455 110.775 97.665 111.295 ;
        RECT 97.835 110.945 99.045 111.465 ;
        RECT 99.675 111.390 99.965 112.555 ;
        RECT 100.135 112.120 105.480 112.555 ;
        RECT 74.375 110.005 79.720 110.550 ;
        RECT 79.895 110.005 85.240 110.550 ;
        RECT 85.415 110.005 90.760 110.550 ;
        RECT 90.935 110.005 96.280 110.550 ;
        RECT 96.455 110.005 99.045 110.775 ;
        RECT 99.675 110.005 99.965 110.730 ;
        RECT 101.720 110.550 102.060 111.380 ;
        RECT 103.540 110.870 103.890 112.120 ;
        RECT 105.655 111.465 107.325 112.555 ;
        RECT 105.655 110.775 106.405 111.295 ;
        RECT 106.575 110.945 107.325 111.465 ;
        RECT 107.955 111.465 109.165 112.555 ;
        RECT 107.955 110.925 108.475 111.465 ;
        RECT 100.135 110.005 105.480 110.550 ;
        RECT 105.655 110.005 107.325 110.775 ;
        RECT 108.645 110.755 109.165 111.295 ;
        RECT 107.955 110.005 109.165 110.755 ;
        RECT 35.190 109.835 109.250 110.005 ;
        RECT 35.275 109.085 36.485 109.835 ;
        RECT 36.655 109.290 42.000 109.835 ;
        RECT 42.175 109.290 47.520 109.835 ;
        RECT 47.695 109.290 53.040 109.835 ;
        RECT 53.215 109.290 58.560 109.835 ;
        RECT 35.275 108.545 35.795 109.085 ;
        RECT 35.965 108.375 36.485 108.915 ;
        RECT 38.240 108.460 38.580 109.290 ;
        RECT 35.275 107.285 36.485 108.375 ;
        RECT 40.060 107.720 40.410 108.970 ;
        RECT 43.760 108.460 44.100 109.290 ;
        RECT 45.580 107.720 45.930 108.970 ;
        RECT 49.280 108.460 49.620 109.290 ;
        RECT 51.100 107.720 51.450 108.970 ;
        RECT 54.800 108.460 55.140 109.290 ;
        RECT 58.735 109.065 60.405 109.835 ;
        RECT 61.035 109.110 61.325 109.835 ;
        RECT 61.495 109.290 66.840 109.835 ;
        RECT 67.015 109.290 72.360 109.835 ;
        RECT 72.535 109.290 77.880 109.835 ;
        RECT 78.055 109.290 83.400 109.835 ;
        RECT 56.620 107.720 56.970 108.970 ;
        RECT 58.735 108.545 59.485 109.065 ;
        RECT 59.655 108.375 60.405 108.895 ;
        RECT 63.080 108.460 63.420 109.290 ;
        RECT 36.655 107.285 42.000 107.720 ;
        RECT 42.175 107.285 47.520 107.720 ;
        RECT 47.695 107.285 53.040 107.720 ;
        RECT 53.215 107.285 58.560 107.720 ;
        RECT 58.735 107.285 60.405 108.375 ;
        RECT 61.035 107.285 61.325 108.450 ;
        RECT 64.900 107.720 65.250 108.970 ;
        RECT 68.600 108.460 68.940 109.290 ;
        RECT 70.420 107.720 70.770 108.970 ;
        RECT 74.120 108.460 74.460 109.290 ;
        RECT 75.940 107.720 76.290 108.970 ;
        RECT 79.640 108.460 79.980 109.290 ;
        RECT 83.575 109.065 86.165 109.835 ;
        RECT 86.795 109.110 87.085 109.835 ;
        RECT 87.255 109.290 92.600 109.835 ;
        RECT 92.775 109.290 98.120 109.835 ;
        RECT 98.295 109.290 103.640 109.835 ;
        RECT 81.460 107.720 81.810 108.970 ;
        RECT 83.575 108.545 84.785 109.065 ;
        RECT 84.955 108.375 86.165 108.895 ;
        RECT 88.840 108.460 89.180 109.290 ;
        RECT 61.495 107.285 66.840 107.720 ;
        RECT 67.015 107.285 72.360 107.720 ;
        RECT 72.535 107.285 77.880 107.720 ;
        RECT 78.055 107.285 83.400 107.720 ;
        RECT 83.575 107.285 86.165 108.375 ;
        RECT 86.795 107.285 87.085 108.450 ;
        RECT 90.660 107.720 91.010 108.970 ;
        RECT 94.360 108.460 94.700 109.290 ;
        RECT 96.180 107.720 96.530 108.970 ;
        RECT 99.880 108.460 100.220 109.290 ;
        RECT 103.815 109.065 107.325 109.835 ;
        RECT 107.955 109.085 109.165 109.835 ;
        RECT 101.700 107.720 102.050 108.970 ;
        RECT 103.815 108.545 105.465 109.065 ;
        RECT 105.635 108.375 107.325 108.895 ;
        RECT 87.255 107.285 92.600 107.720 ;
        RECT 92.775 107.285 98.120 107.720 ;
        RECT 98.295 107.285 103.640 107.720 ;
        RECT 103.815 107.285 107.325 108.375 ;
        RECT 107.955 108.375 108.475 108.915 ;
        RECT 108.645 108.545 109.165 109.085 ;
        RECT 107.955 107.285 109.165 108.375 ;
        RECT 35.190 107.115 109.250 107.285 ;
        RECT 35.275 106.025 36.485 107.115 ;
        RECT 36.655 106.680 42.000 107.115 ;
        RECT 42.175 106.680 47.520 107.115 ;
        RECT 35.275 105.315 35.795 105.855 ;
        RECT 35.965 105.485 36.485 106.025 ;
        RECT 35.275 104.565 36.485 105.315 ;
        RECT 38.240 105.110 38.580 105.940 ;
        RECT 40.060 105.430 40.410 106.680 ;
        RECT 43.760 105.110 44.100 105.940 ;
        RECT 45.580 105.430 45.930 106.680 ;
        RECT 48.155 105.950 48.445 107.115 ;
        RECT 48.615 106.680 53.960 107.115 ;
        RECT 54.135 106.680 59.480 107.115 ;
        RECT 59.655 106.680 65.000 107.115 ;
        RECT 65.175 106.680 70.520 107.115 ;
        RECT 36.655 104.565 42.000 105.110 ;
        RECT 42.175 104.565 47.520 105.110 ;
        RECT 48.155 104.565 48.445 105.290 ;
        RECT 50.200 105.110 50.540 105.940 ;
        RECT 52.020 105.430 52.370 106.680 ;
        RECT 55.720 105.110 56.060 105.940 ;
        RECT 57.540 105.430 57.890 106.680 ;
        RECT 61.240 105.110 61.580 105.940 ;
        RECT 63.060 105.430 63.410 106.680 ;
        RECT 66.760 105.110 67.100 105.940 ;
        RECT 68.580 105.430 68.930 106.680 ;
        RECT 70.695 106.025 73.285 107.115 ;
        RECT 70.695 105.335 71.905 105.855 ;
        RECT 72.075 105.505 73.285 106.025 ;
        RECT 73.915 105.950 74.205 107.115 ;
        RECT 74.375 106.680 79.720 107.115 ;
        RECT 79.895 106.680 85.240 107.115 ;
        RECT 85.415 106.680 90.760 107.115 ;
        RECT 90.935 106.680 96.280 107.115 ;
        RECT 48.615 104.565 53.960 105.110 ;
        RECT 54.135 104.565 59.480 105.110 ;
        RECT 59.655 104.565 65.000 105.110 ;
        RECT 65.175 104.565 70.520 105.110 ;
        RECT 70.695 104.565 73.285 105.335 ;
        RECT 73.915 104.565 74.205 105.290 ;
        RECT 75.960 105.110 76.300 105.940 ;
        RECT 77.780 105.430 78.130 106.680 ;
        RECT 81.480 105.110 81.820 105.940 ;
        RECT 83.300 105.430 83.650 106.680 ;
        RECT 87.000 105.110 87.340 105.940 ;
        RECT 88.820 105.430 89.170 106.680 ;
        RECT 92.520 105.110 92.860 105.940 ;
        RECT 94.340 105.430 94.690 106.680 ;
        RECT 96.455 106.025 99.045 107.115 ;
        RECT 96.455 105.335 97.665 105.855 ;
        RECT 97.835 105.505 99.045 106.025 ;
        RECT 99.675 105.950 99.965 107.115 ;
        RECT 100.135 106.680 105.480 107.115 ;
        RECT 74.375 104.565 79.720 105.110 ;
        RECT 79.895 104.565 85.240 105.110 ;
        RECT 85.415 104.565 90.760 105.110 ;
        RECT 90.935 104.565 96.280 105.110 ;
        RECT 96.455 104.565 99.045 105.335 ;
        RECT 99.675 104.565 99.965 105.290 ;
        RECT 101.720 105.110 102.060 105.940 ;
        RECT 103.540 105.430 103.890 106.680 ;
        RECT 105.655 106.025 107.325 107.115 ;
        RECT 105.655 105.335 106.405 105.855 ;
        RECT 106.575 105.505 107.325 106.025 ;
        RECT 107.955 106.025 109.165 107.115 ;
        RECT 107.955 105.485 108.475 106.025 ;
        RECT 100.135 104.565 105.480 105.110 ;
        RECT 105.655 104.565 107.325 105.335 ;
        RECT 108.645 105.315 109.165 105.855 ;
        RECT 107.955 104.565 109.165 105.315 ;
        RECT 35.190 104.395 109.250 104.565 ;
        RECT 35.275 103.645 36.485 104.395 ;
        RECT 36.655 103.850 42.000 104.395 ;
        RECT 42.175 103.850 47.520 104.395 ;
        RECT 47.695 103.850 53.040 104.395 ;
        RECT 53.215 103.850 58.560 104.395 ;
        RECT 35.275 103.105 35.795 103.645 ;
        RECT 35.965 102.935 36.485 103.475 ;
        RECT 38.240 103.020 38.580 103.850 ;
        RECT 35.275 101.845 36.485 102.935 ;
        RECT 40.060 102.280 40.410 103.530 ;
        RECT 43.760 103.020 44.100 103.850 ;
        RECT 45.580 102.280 45.930 103.530 ;
        RECT 49.280 103.020 49.620 103.850 ;
        RECT 51.100 102.280 51.450 103.530 ;
        RECT 54.800 103.020 55.140 103.850 ;
        RECT 58.735 103.625 60.405 104.395 ;
        RECT 61.035 103.670 61.325 104.395 ;
        RECT 61.495 103.850 66.840 104.395 ;
        RECT 67.015 103.850 72.360 104.395 ;
        RECT 72.535 103.850 77.880 104.395 ;
        RECT 78.055 103.850 83.400 104.395 ;
        RECT 56.620 102.280 56.970 103.530 ;
        RECT 58.735 103.105 59.485 103.625 ;
        RECT 59.655 102.935 60.405 103.455 ;
        RECT 63.080 103.020 63.420 103.850 ;
        RECT 36.655 101.845 42.000 102.280 ;
        RECT 42.175 101.845 47.520 102.280 ;
        RECT 47.695 101.845 53.040 102.280 ;
        RECT 53.215 101.845 58.560 102.280 ;
        RECT 58.735 101.845 60.405 102.935 ;
        RECT 61.035 101.845 61.325 103.010 ;
        RECT 64.900 102.280 65.250 103.530 ;
        RECT 68.600 103.020 68.940 103.850 ;
        RECT 70.420 102.280 70.770 103.530 ;
        RECT 74.120 103.020 74.460 103.850 ;
        RECT 75.940 102.280 76.290 103.530 ;
        RECT 79.640 103.020 79.980 103.850 ;
        RECT 83.575 103.625 86.165 104.395 ;
        RECT 86.795 103.670 87.085 104.395 ;
        RECT 87.255 103.850 92.600 104.395 ;
        RECT 92.775 103.850 98.120 104.395 ;
        RECT 98.295 103.850 103.640 104.395 ;
        RECT 81.460 102.280 81.810 103.530 ;
        RECT 83.575 103.105 84.785 103.625 ;
        RECT 84.955 102.935 86.165 103.455 ;
        RECT 88.840 103.020 89.180 103.850 ;
        RECT 61.495 101.845 66.840 102.280 ;
        RECT 67.015 101.845 72.360 102.280 ;
        RECT 72.535 101.845 77.880 102.280 ;
        RECT 78.055 101.845 83.400 102.280 ;
        RECT 83.575 101.845 86.165 102.935 ;
        RECT 86.795 101.845 87.085 103.010 ;
        RECT 90.660 102.280 91.010 103.530 ;
        RECT 94.360 103.020 94.700 103.850 ;
        RECT 96.180 102.280 96.530 103.530 ;
        RECT 99.880 103.020 100.220 103.850 ;
        RECT 103.815 103.625 107.325 104.395 ;
        RECT 107.955 103.645 109.165 104.395 ;
        RECT 101.700 102.280 102.050 103.530 ;
        RECT 103.815 103.105 105.465 103.625 ;
        RECT 105.635 102.935 107.325 103.455 ;
        RECT 87.255 101.845 92.600 102.280 ;
        RECT 92.775 101.845 98.120 102.280 ;
        RECT 98.295 101.845 103.640 102.280 ;
        RECT 103.815 101.845 107.325 102.935 ;
        RECT 107.955 102.935 108.475 103.475 ;
        RECT 108.645 103.105 109.165 103.645 ;
        RECT 107.955 101.845 109.165 102.935 ;
        RECT 35.190 101.675 109.250 101.845 ;
        RECT 35.275 100.585 36.485 101.675 ;
        RECT 36.655 101.240 42.000 101.675 ;
        RECT 42.175 101.240 47.520 101.675 ;
        RECT 35.275 99.875 35.795 100.415 ;
        RECT 35.965 100.045 36.485 100.585 ;
        RECT 35.275 99.125 36.485 99.875 ;
        RECT 38.240 99.670 38.580 100.500 ;
        RECT 40.060 99.990 40.410 101.240 ;
        RECT 43.760 99.670 44.100 100.500 ;
        RECT 45.580 99.990 45.930 101.240 ;
        RECT 48.155 100.510 48.445 101.675 ;
        RECT 48.615 101.240 53.960 101.675 ;
        RECT 54.135 101.240 59.480 101.675 ;
        RECT 59.655 101.240 65.000 101.675 ;
        RECT 65.175 101.240 70.520 101.675 ;
        RECT 36.655 99.125 42.000 99.670 ;
        RECT 42.175 99.125 47.520 99.670 ;
        RECT 48.155 99.125 48.445 99.850 ;
        RECT 50.200 99.670 50.540 100.500 ;
        RECT 52.020 99.990 52.370 101.240 ;
        RECT 55.720 99.670 56.060 100.500 ;
        RECT 57.540 99.990 57.890 101.240 ;
        RECT 61.240 99.670 61.580 100.500 ;
        RECT 63.060 99.990 63.410 101.240 ;
        RECT 66.760 99.670 67.100 100.500 ;
        RECT 68.580 99.990 68.930 101.240 ;
        RECT 70.695 100.585 73.285 101.675 ;
        RECT 70.695 99.895 71.905 100.415 ;
        RECT 72.075 100.065 73.285 100.585 ;
        RECT 73.915 100.510 74.205 101.675 ;
        RECT 74.375 101.240 79.720 101.675 ;
        RECT 79.895 101.240 85.240 101.675 ;
        RECT 85.415 101.240 90.760 101.675 ;
        RECT 90.935 101.240 96.280 101.675 ;
        RECT 48.615 99.125 53.960 99.670 ;
        RECT 54.135 99.125 59.480 99.670 ;
        RECT 59.655 99.125 65.000 99.670 ;
        RECT 65.175 99.125 70.520 99.670 ;
        RECT 70.695 99.125 73.285 99.895 ;
        RECT 73.915 99.125 74.205 99.850 ;
        RECT 75.960 99.670 76.300 100.500 ;
        RECT 77.780 99.990 78.130 101.240 ;
        RECT 81.480 99.670 81.820 100.500 ;
        RECT 83.300 99.990 83.650 101.240 ;
        RECT 87.000 99.670 87.340 100.500 ;
        RECT 88.820 99.990 89.170 101.240 ;
        RECT 92.520 99.670 92.860 100.500 ;
        RECT 94.340 99.990 94.690 101.240 ;
        RECT 96.455 100.585 99.045 101.675 ;
        RECT 96.455 99.895 97.665 100.415 ;
        RECT 97.835 100.065 99.045 100.585 ;
        RECT 99.675 100.510 99.965 101.675 ;
        RECT 100.135 101.240 105.480 101.675 ;
        RECT 74.375 99.125 79.720 99.670 ;
        RECT 79.895 99.125 85.240 99.670 ;
        RECT 85.415 99.125 90.760 99.670 ;
        RECT 90.935 99.125 96.280 99.670 ;
        RECT 96.455 99.125 99.045 99.895 ;
        RECT 99.675 99.125 99.965 99.850 ;
        RECT 101.720 99.670 102.060 100.500 ;
        RECT 103.540 99.990 103.890 101.240 ;
        RECT 105.655 100.585 107.325 101.675 ;
        RECT 105.655 99.895 106.405 100.415 ;
        RECT 106.575 100.065 107.325 100.585 ;
        RECT 107.955 100.585 109.165 101.675 ;
        RECT 107.955 100.045 108.475 100.585 ;
        RECT 100.135 99.125 105.480 99.670 ;
        RECT 105.655 99.125 107.325 99.895 ;
        RECT 108.645 99.875 109.165 100.415 ;
        RECT 107.955 99.125 109.165 99.875 ;
        RECT 35.190 98.955 109.250 99.125 ;
        RECT 35.275 98.205 36.485 98.955 ;
        RECT 36.655 98.410 42.000 98.955 ;
        RECT 42.175 98.410 47.520 98.955 ;
        RECT 47.695 98.410 53.040 98.955 ;
        RECT 53.215 98.410 58.560 98.955 ;
        RECT 35.275 97.665 35.795 98.205 ;
        RECT 35.965 97.495 36.485 98.035 ;
        RECT 38.240 97.580 38.580 98.410 ;
        RECT 35.275 96.405 36.485 97.495 ;
        RECT 40.060 96.840 40.410 98.090 ;
        RECT 43.760 97.580 44.100 98.410 ;
        RECT 45.580 96.840 45.930 98.090 ;
        RECT 49.280 97.580 49.620 98.410 ;
        RECT 51.100 96.840 51.450 98.090 ;
        RECT 54.800 97.580 55.140 98.410 ;
        RECT 58.735 98.185 60.405 98.955 ;
        RECT 61.035 98.230 61.325 98.955 ;
        RECT 61.495 98.410 66.840 98.955 ;
        RECT 67.015 98.410 72.360 98.955 ;
        RECT 72.535 98.410 77.880 98.955 ;
        RECT 78.055 98.410 83.400 98.955 ;
        RECT 56.620 96.840 56.970 98.090 ;
        RECT 58.735 97.665 59.485 98.185 ;
        RECT 59.655 97.495 60.405 98.015 ;
        RECT 63.080 97.580 63.420 98.410 ;
        RECT 36.655 96.405 42.000 96.840 ;
        RECT 42.175 96.405 47.520 96.840 ;
        RECT 47.695 96.405 53.040 96.840 ;
        RECT 53.215 96.405 58.560 96.840 ;
        RECT 58.735 96.405 60.405 97.495 ;
        RECT 61.035 96.405 61.325 97.570 ;
        RECT 64.900 96.840 65.250 98.090 ;
        RECT 68.600 97.580 68.940 98.410 ;
        RECT 70.420 96.840 70.770 98.090 ;
        RECT 74.120 97.580 74.460 98.410 ;
        RECT 75.940 96.840 76.290 98.090 ;
        RECT 79.640 97.580 79.980 98.410 ;
        RECT 83.575 98.185 86.165 98.955 ;
        RECT 86.795 98.230 87.085 98.955 ;
        RECT 87.255 98.410 92.600 98.955 ;
        RECT 92.775 98.410 98.120 98.955 ;
        RECT 98.295 98.410 103.640 98.955 ;
        RECT 81.460 96.840 81.810 98.090 ;
        RECT 83.575 97.665 84.785 98.185 ;
        RECT 84.955 97.495 86.165 98.015 ;
        RECT 88.840 97.580 89.180 98.410 ;
        RECT 61.495 96.405 66.840 96.840 ;
        RECT 67.015 96.405 72.360 96.840 ;
        RECT 72.535 96.405 77.880 96.840 ;
        RECT 78.055 96.405 83.400 96.840 ;
        RECT 83.575 96.405 86.165 97.495 ;
        RECT 86.795 96.405 87.085 97.570 ;
        RECT 90.660 96.840 91.010 98.090 ;
        RECT 94.360 97.580 94.700 98.410 ;
        RECT 96.180 96.840 96.530 98.090 ;
        RECT 99.880 97.580 100.220 98.410 ;
        RECT 103.815 98.185 107.325 98.955 ;
        RECT 107.955 98.205 109.165 98.955 ;
        RECT 101.700 96.840 102.050 98.090 ;
        RECT 103.815 97.665 105.465 98.185 ;
        RECT 105.635 97.495 107.325 98.015 ;
        RECT 87.255 96.405 92.600 96.840 ;
        RECT 92.775 96.405 98.120 96.840 ;
        RECT 98.295 96.405 103.640 96.840 ;
        RECT 103.815 96.405 107.325 97.495 ;
        RECT 107.955 97.495 108.475 98.035 ;
        RECT 108.645 97.665 109.165 98.205 ;
        RECT 107.955 96.405 109.165 97.495 ;
        RECT 35.190 96.235 109.250 96.405 ;
        RECT 35.275 95.145 36.485 96.235 ;
        RECT 36.655 95.800 42.000 96.235 ;
        RECT 42.175 95.800 47.520 96.235 ;
        RECT 35.275 94.435 35.795 94.975 ;
        RECT 35.965 94.605 36.485 95.145 ;
        RECT 35.275 93.685 36.485 94.435 ;
        RECT 38.240 94.230 38.580 95.060 ;
        RECT 40.060 94.550 40.410 95.800 ;
        RECT 43.760 94.230 44.100 95.060 ;
        RECT 45.580 94.550 45.930 95.800 ;
        RECT 48.155 95.070 48.445 96.235 ;
        RECT 48.615 95.800 53.960 96.235 ;
        RECT 54.135 95.800 59.480 96.235 ;
        RECT 59.655 95.800 65.000 96.235 ;
        RECT 65.175 95.800 70.520 96.235 ;
        RECT 36.655 93.685 42.000 94.230 ;
        RECT 42.175 93.685 47.520 94.230 ;
        RECT 48.155 93.685 48.445 94.410 ;
        RECT 50.200 94.230 50.540 95.060 ;
        RECT 52.020 94.550 52.370 95.800 ;
        RECT 55.720 94.230 56.060 95.060 ;
        RECT 57.540 94.550 57.890 95.800 ;
        RECT 61.240 94.230 61.580 95.060 ;
        RECT 63.060 94.550 63.410 95.800 ;
        RECT 66.760 94.230 67.100 95.060 ;
        RECT 68.580 94.550 68.930 95.800 ;
        RECT 70.695 95.145 73.285 96.235 ;
        RECT 70.695 94.455 71.905 94.975 ;
        RECT 72.075 94.625 73.285 95.145 ;
        RECT 73.915 95.070 74.205 96.235 ;
        RECT 74.375 95.800 79.720 96.235 ;
        RECT 79.895 95.800 85.240 96.235 ;
        RECT 85.415 95.800 90.760 96.235 ;
        RECT 90.935 95.800 96.280 96.235 ;
        RECT 48.615 93.685 53.960 94.230 ;
        RECT 54.135 93.685 59.480 94.230 ;
        RECT 59.655 93.685 65.000 94.230 ;
        RECT 65.175 93.685 70.520 94.230 ;
        RECT 70.695 93.685 73.285 94.455 ;
        RECT 73.915 93.685 74.205 94.410 ;
        RECT 75.960 94.230 76.300 95.060 ;
        RECT 77.780 94.550 78.130 95.800 ;
        RECT 81.480 94.230 81.820 95.060 ;
        RECT 83.300 94.550 83.650 95.800 ;
        RECT 87.000 94.230 87.340 95.060 ;
        RECT 88.820 94.550 89.170 95.800 ;
        RECT 92.520 94.230 92.860 95.060 ;
        RECT 94.340 94.550 94.690 95.800 ;
        RECT 96.455 95.145 99.045 96.235 ;
        RECT 96.455 94.455 97.665 94.975 ;
        RECT 97.835 94.625 99.045 95.145 ;
        RECT 99.675 95.070 99.965 96.235 ;
        RECT 100.135 95.800 105.480 96.235 ;
        RECT 74.375 93.685 79.720 94.230 ;
        RECT 79.895 93.685 85.240 94.230 ;
        RECT 85.415 93.685 90.760 94.230 ;
        RECT 90.935 93.685 96.280 94.230 ;
        RECT 96.455 93.685 99.045 94.455 ;
        RECT 99.675 93.685 99.965 94.410 ;
        RECT 101.720 94.230 102.060 95.060 ;
        RECT 103.540 94.550 103.890 95.800 ;
        RECT 105.655 95.145 107.325 96.235 ;
        RECT 105.655 94.455 106.405 94.975 ;
        RECT 106.575 94.625 107.325 95.145 ;
        RECT 107.955 95.145 109.165 96.235 ;
        RECT 107.955 94.605 108.475 95.145 ;
        RECT 100.135 93.685 105.480 94.230 ;
        RECT 105.655 93.685 107.325 94.455 ;
        RECT 108.645 94.435 109.165 94.975 ;
        RECT 107.955 93.685 109.165 94.435 ;
        RECT 35.190 93.515 109.250 93.685 ;
        RECT 35.275 92.765 36.485 93.515 ;
        RECT 36.655 92.970 42.000 93.515 ;
        RECT 42.175 92.970 47.520 93.515 ;
        RECT 47.695 92.970 53.040 93.515 ;
        RECT 53.215 92.970 58.560 93.515 ;
        RECT 35.275 92.225 35.795 92.765 ;
        RECT 35.965 92.055 36.485 92.595 ;
        RECT 38.240 92.140 38.580 92.970 ;
        RECT 35.275 90.965 36.485 92.055 ;
        RECT 40.060 91.400 40.410 92.650 ;
        RECT 43.760 92.140 44.100 92.970 ;
        RECT 45.580 91.400 45.930 92.650 ;
        RECT 49.280 92.140 49.620 92.970 ;
        RECT 51.100 91.400 51.450 92.650 ;
        RECT 54.800 92.140 55.140 92.970 ;
        RECT 58.735 92.745 60.405 93.515 ;
        RECT 61.035 92.790 61.325 93.515 ;
        RECT 61.495 92.970 66.840 93.515 ;
        RECT 67.015 92.970 72.360 93.515 ;
        RECT 72.535 92.970 77.880 93.515 ;
        RECT 78.055 92.970 83.400 93.515 ;
        RECT 56.620 91.400 56.970 92.650 ;
        RECT 58.735 92.225 59.485 92.745 ;
        RECT 59.655 92.055 60.405 92.575 ;
        RECT 63.080 92.140 63.420 92.970 ;
        RECT 36.655 90.965 42.000 91.400 ;
        RECT 42.175 90.965 47.520 91.400 ;
        RECT 47.695 90.965 53.040 91.400 ;
        RECT 53.215 90.965 58.560 91.400 ;
        RECT 58.735 90.965 60.405 92.055 ;
        RECT 61.035 90.965 61.325 92.130 ;
        RECT 64.900 91.400 65.250 92.650 ;
        RECT 68.600 92.140 68.940 92.970 ;
        RECT 70.420 91.400 70.770 92.650 ;
        RECT 74.120 92.140 74.460 92.970 ;
        RECT 75.940 91.400 76.290 92.650 ;
        RECT 79.640 92.140 79.980 92.970 ;
        RECT 83.575 92.745 86.165 93.515 ;
        RECT 86.795 92.790 87.085 93.515 ;
        RECT 87.255 92.970 92.600 93.515 ;
        RECT 92.775 92.970 98.120 93.515 ;
        RECT 98.295 92.970 103.640 93.515 ;
        RECT 81.460 91.400 81.810 92.650 ;
        RECT 83.575 92.225 84.785 92.745 ;
        RECT 84.955 92.055 86.165 92.575 ;
        RECT 88.840 92.140 89.180 92.970 ;
        RECT 61.495 90.965 66.840 91.400 ;
        RECT 67.015 90.965 72.360 91.400 ;
        RECT 72.535 90.965 77.880 91.400 ;
        RECT 78.055 90.965 83.400 91.400 ;
        RECT 83.575 90.965 86.165 92.055 ;
        RECT 86.795 90.965 87.085 92.130 ;
        RECT 90.660 91.400 91.010 92.650 ;
        RECT 94.360 92.140 94.700 92.970 ;
        RECT 96.180 91.400 96.530 92.650 ;
        RECT 99.880 92.140 100.220 92.970 ;
        RECT 103.815 92.745 107.325 93.515 ;
        RECT 107.955 92.765 109.165 93.515 ;
        RECT 101.700 91.400 102.050 92.650 ;
        RECT 103.815 92.225 105.465 92.745 ;
        RECT 105.635 92.055 107.325 92.575 ;
        RECT 87.255 90.965 92.600 91.400 ;
        RECT 92.775 90.965 98.120 91.400 ;
        RECT 98.295 90.965 103.640 91.400 ;
        RECT 103.815 90.965 107.325 92.055 ;
        RECT 107.955 92.055 108.475 92.595 ;
        RECT 108.645 92.225 109.165 92.765 ;
        RECT 107.955 90.965 109.165 92.055 ;
        RECT 35.190 90.795 109.250 90.965 ;
        RECT 35.275 89.705 36.485 90.795 ;
        RECT 36.655 90.360 42.000 90.795 ;
        RECT 42.175 90.360 47.520 90.795 ;
        RECT 35.275 88.995 35.795 89.535 ;
        RECT 35.965 89.165 36.485 89.705 ;
        RECT 35.275 88.245 36.485 88.995 ;
        RECT 38.240 88.790 38.580 89.620 ;
        RECT 40.060 89.110 40.410 90.360 ;
        RECT 43.760 88.790 44.100 89.620 ;
        RECT 45.580 89.110 45.930 90.360 ;
        RECT 48.155 89.630 48.445 90.795 ;
        RECT 48.615 90.360 53.960 90.795 ;
        RECT 54.135 90.360 59.480 90.795 ;
        RECT 59.655 90.360 65.000 90.795 ;
        RECT 65.175 90.360 70.520 90.795 ;
        RECT 36.655 88.245 42.000 88.790 ;
        RECT 42.175 88.245 47.520 88.790 ;
        RECT 48.155 88.245 48.445 88.970 ;
        RECT 50.200 88.790 50.540 89.620 ;
        RECT 52.020 89.110 52.370 90.360 ;
        RECT 55.720 88.790 56.060 89.620 ;
        RECT 57.540 89.110 57.890 90.360 ;
        RECT 61.240 88.790 61.580 89.620 ;
        RECT 63.060 89.110 63.410 90.360 ;
        RECT 66.760 88.790 67.100 89.620 ;
        RECT 68.580 89.110 68.930 90.360 ;
        RECT 70.695 89.705 73.285 90.795 ;
        RECT 70.695 89.015 71.905 89.535 ;
        RECT 72.075 89.185 73.285 89.705 ;
        RECT 73.915 89.630 74.205 90.795 ;
        RECT 74.375 90.360 79.720 90.795 ;
        RECT 79.895 90.360 85.240 90.795 ;
        RECT 85.415 90.360 90.760 90.795 ;
        RECT 90.935 90.360 96.280 90.795 ;
        RECT 48.615 88.245 53.960 88.790 ;
        RECT 54.135 88.245 59.480 88.790 ;
        RECT 59.655 88.245 65.000 88.790 ;
        RECT 65.175 88.245 70.520 88.790 ;
        RECT 70.695 88.245 73.285 89.015 ;
        RECT 73.915 88.245 74.205 88.970 ;
        RECT 75.960 88.790 76.300 89.620 ;
        RECT 77.780 89.110 78.130 90.360 ;
        RECT 81.480 88.790 81.820 89.620 ;
        RECT 83.300 89.110 83.650 90.360 ;
        RECT 87.000 88.790 87.340 89.620 ;
        RECT 88.820 89.110 89.170 90.360 ;
        RECT 92.520 88.790 92.860 89.620 ;
        RECT 94.340 89.110 94.690 90.360 ;
        RECT 96.455 89.705 99.045 90.795 ;
        RECT 96.455 89.015 97.665 89.535 ;
        RECT 97.835 89.185 99.045 89.705 ;
        RECT 99.675 89.630 99.965 90.795 ;
        RECT 100.135 90.360 105.480 90.795 ;
        RECT 74.375 88.245 79.720 88.790 ;
        RECT 79.895 88.245 85.240 88.790 ;
        RECT 85.415 88.245 90.760 88.790 ;
        RECT 90.935 88.245 96.280 88.790 ;
        RECT 96.455 88.245 99.045 89.015 ;
        RECT 99.675 88.245 99.965 88.970 ;
        RECT 101.720 88.790 102.060 89.620 ;
        RECT 103.540 89.110 103.890 90.360 ;
        RECT 105.655 89.705 107.325 90.795 ;
        RECT 105.655 89.015 106.405 89.535 ;
        RECT 106.575 89.185 107.325 89.705 ;
        RECT 107.955 89.705 109.165 90.795 ;
        RECT 107.955 89.165 108.475 89.705 ;
        RECT 100.135 88.245 105.480 88.790 ;
        RECT 105.655 88.245 107.325 89.015 ;
        RECT 108.645 88.995 109.165 89.535 ;
        RECT 107.955 88.245 109.165 88.995 ;
        RECT 35.190 88.075 109.250 88.245 ;
        RECT 35.275 87.325 36.485 88.075 ;
        RECT 36.655 87.530 42.000 88.075 ;
        RECT 42.175 87.530 47.520 88.075 ;
        RECT 47.695 87.530 53.040 88.075 ;
        RECT 53.215 87.530 58.560 88.075 ;
        RECT 35.275 86.785 35.795 87.325 ;
        RECT 35.965 86.615 36.485 87.155 ;
        RECT 38.240 86.700 38.580 87.530 ;
        RECT 35.275 85.525 36.485 86.615 ;
        RECT 40.060 85.960 40.410 87.210 ;
        RECT 43.760 86.700 44.100 87.530 ;
        RECT 45.580 85.960 45.930 87.210 ;
        RECT 49.280 86.700 49.620 87.530 ;
        RECT 51.100 85.960 51.450 87.210 ;
        RECT 54.800 86.700 55.140 87.530 ;
        RECT 58.735 87.305 60.405 88.075 ;
        RECT 61.035 87.350 61.325 88.075 ;
        RECT 61.495 87.530 66.840 88.075 ;
        RECT 67.015 87.530 72.360 88.075 ;
        RECT 72.535 87.530 77.880 88.075 ;
        RECT 78.055 87.530 83.400 88.075 ;
        RECT 56.620 85.960 56.970 87.210 ;
        RECT 58.735 86.785 59.485 87.305 ;
        RECT 59.655 86.615 60.405 87.135 ;
        RECT 63.080 86.700 63.420 87.530 ;
        RECT 36.655 85.525 42.000 85.960 ;
        RECT 42.175 85.525 47.520 85.960 ;
        RECT 47.695 85.525 53.040 85.960 ;
        RECT 53.215 85.525 58.560 85.960 ;
        RECT 58.735 85.525 60.405 86.615 ;
        RECT 61.035 85.525 61.325 86.690 ;
        RECT 64.900 85.960 65.250 87.210 ;
        RECT 68.600 86.700 68.940 87.530 ;
        RECT 70.420 85.960 70.770 87.210 ;
        RECT 74.120 86.700 74.460 87.530 ;
        RECT 75.940 85.960 76.290 87.210 ;
        RECT 79.640 86.700 79.980 87.530 ;
        RECT 83.575 87.305 86.165 88.075 ;
        RECT 86.795 87.350 87.085 88.075 ;
        RECT 87.255 87.530 92.600 88.075 ;
        RECT 92.775 87.530 98.120 88.075 ;
        RECT 98.295 87.530 103.640 88.075 ;
        RECT 81.460 85.960 81.810 87.210 ;
        RECT 83.575 86.785 84.785 87.305 ;
        RECT 84.955 86.615 86.165 87.135 ;
        RECT 88.840 86.700 89.180 87.530 ;
        RECT 61.495 85.525 66.840 85.960 ;
        RECT 67.015 85.525 72.360 85.960 ;
        RECT 72.535 85.525 77.880 85.960 ;
        RECT 78.055 85.525 83.400 85.960 ;
        RECT 83.575 85.525 86.165 86.615 ;
        RECT 86.795 85.525 87.085 86.690 ;
        RECT 90.660 85.960 91.010 87.210 ;
        RECT 94.360 86.700 94.700 87.530 ;
        RECT 96.180 85.960 96.530 87.210 ;
        RECT 99.880 86.700 100.220 87.530 ;
        RECT 103.815 87.305 107.325 88.075 ;
        RECT 107.955 87.325 109.165 88.075 ;
        RECT 101.700 85.960 102.050 87.210 ;
        RECT 103.815 86.785 105.465 87.305 ;
        RECT 105.635 86.615 107.325 87.135 ;
        RECT 87.255 85.525 92.600 85.960 ;
        RECT 92.775 85.525 98.120 85.960 ;
        RECT 98.295 85.525 103.640 85.960 ;
        RECT 103.815 85.525 107.325 86.615 ;
        RECT 107.955 86.615 108.475 87.155 ;
        RECT 108.645 86.785 109.165 87.325 ;
        RECT 107.955 85.525 109.165 86.615 ;
        RECT 35.190 85.355 109.250 85.525 ;
        RECT 35.275 84.265 36.485 85.355 ;
        RECT 36.655 84.920 42.000 85.355 ;
        RECT 42.175 84.920 47.520 85.355 ;
        RECT 35.275 83.555 35.795 84.095 ;
        RECT 35.965 83.725 36.485 84.265 ;
        RECT 35.275 82.805 36.485 83.555 ;
        RECT 38.240 83.350 38.580 84.180 ;
        RECT 40.060 83.670 40.410 84.920 ;
        RECT 43.760 83.350 44.100 84.180 ;
        RECT 45.580 83.670 45.930 84.920 ;
        RECT 48.155 84.190 48.445 85.355 ;
        RECT 48.615 84.920 53.960 85.355 ;
        RECT 54.135 84.920 59.480 85.355 ;
        RECT 36.655 82.805 42.000 83.350 ;
        RECT 42.175 82.805 47.520 83.350 ;
        RECT 48.155 82.805 48.445 83.530 ;
        RECT 50.200 83.350 50.540 84.180 ;
        RECT 52.020 83.670 52.370 84.920 ;
        RECT 55.720 83.350 56.060 84.180 ;
        RECT 57.540 83.670 57.890 84.920 ;
        RECT 59.655 84.265 60.865 85.355 ;
        RECT 59.655 83.555 60.175 84.095 ;
        RECT 60.345 83.725 60.865 84.265 ;
        RECT 61.035 84.190 61.325 85.355 ;
        RECT 61.495 84.920 66.840 85.355 ;
        RECT 67.015 84.920 72.360 85.355 ;
        RECT 48.615 82.805 53.960 83.350 ;
        RECT 54.135 82.805 59.480 83.350 ;
        RECT 59.655 82.805 60.865 83.555 ;
        RECT 61.035 82.805 61.325 83.530 ;
        RECT 63.080 83.350 63.420 84.180 ;
        RECT 64.900 83.670 65.250 84.920 ;
        RECT 68.600 83.350 68.940 84.180 ;
        RECT 70.420 83.670 70.770 84.920 ;
        RECT 72.535 84.265 73.745 85.355 ;
        RECT 72.535 83.555 73.055 84.095 ;
        RECT 73.225 83.725 73.745 84.265 ;
        RECT 73.915 84.190 74.205 85.355 ;
        RECT 74.375 84.385 74.645 85.155 ;
        RECT 74.815 84.575 75.145 85.355 ;
        RECT 75.350 84.750 75.535 85.155 ;
        RECT 75.705 84.930 76.040 85.355 ;
        RECT 76.215 84.920 81.560 85.355 ;
        RECT 75.350 84.575 76.015 84.750 ;
        RECT 74.375 84.215 75.505 84.385 ;
        RECT 61.495 82.805 66.840 83.350 ;
        RECT 67.015 82.805 72.360 83.350 ;
        RECT 72.535 82.805 73.745 83.555 ;
        RECT 73.915 82.805 74.205 83.530 ;
        RECT 74.375 83.305 74.545 84.215 ;
        RECT 74.715 83.465 75.075 84.045 ;
        RECT 75.255 83.715 75.505 84.215 ;
        RECT 75.675 83.545 76.015 84.575 ;
        RECT 75.330 83.375 76.015 83.545 ;
        RECT 74.375 82.975 74.635 83.305 ;
        RECT 74.845 82.805 75.120 83.285 ;
        RECT 75.330 82.975 75.535 83.375 ;
        RECT 77.800 83.350 78.140 84.180 ;
        RECT 79.620 83.670 79.970 84.920 ;
        RECT 81.735 84.265 85.245 85.355 ;
        RECT 85.415 84.265 86.625 85.355 ;
        RECT 81.735 83.575 83.385 84.095 ;
        RECT 83.555 83.745 85.245 84.265 ;
        RECT 75.705 82.805 76.040 83.205 ;
        RECT 76.215 82.805 81.560 83.350 ;
        RECT 81.735 82.805 85.245 83.575 ;
        RECT 85.415 83.555 85.935 84.095 ;
        RECT 86.105 83.725 86.625 84.265 ;
        RECT 86.795 84.190 87.085 85.355 ;
        RECT 87.255 84.920 92.600 85.355 ;
        RECT 92.775 84.920 98.120 85.355 ;
        RECT 85.415 82.805 86.625 83.555 ;
        RECT 86.795 82.805 87.085 83.530 ;
        RECT 88.840 83.350 89.180 84.180 ;
        RECT 90.660 83.670 91.010 84.920 ;
        RECT 94.360 83.350 94.700 84.180 ;
        RECT 96.180 83.670 96.530 84.920 ;
        RECT 98.295 84.265 99.505 85.355 ;
        RECT 98.295 83.555 98.815 84.095 ;
        RECT 98.985 83.725 99.505 84.265 ;
        RECT 99.675 84.190 99.965 85.355 ;
        RECT 100.135 84.920 105.480 85.355 ;
        RECT 87.255 82.805 92.600 83.350 ;
        RECT 92.775 82.805 98.120 83.350 ;
        RECT 98.295 82.805 99.505 83.555 ;
        RECT 99.675 82.805 99.965 83.530 ;
        RECT 101.720 83.350 102.060 84.180 ;
        RECT 103.540 83.670 103.890 84.920 ;
        RECT 105.655 84.265 107.325 85.355 ;
        RECT 105.655 83.575 106.405 84.095 ;
        RECT 106.575 83.745 107.325 84.265 ;
        RECT 107.955 84.265 109.165 85.355 ;
        RECT 107.955 83.725 108.475 84.265 ;
        RECT 100.135 82.805 105.480 83.350 ;
        RECT 105.655 82.805 107.325 83.575 ;
        RECT 108.645 83.555 109.165 84.095 ;
        RECT 107.955 82.805 109.165 83.555 ;
        RECT 35.190 82.635 109.250 82.805 ;
        RECT 107.140 77.360 110.220 77.530 ;
        RECT 110.840 77.370 113.920 77.540 ;
        RECT 114.550 77.370 117.630 77.540 ;
        RECT 118.260 77.370 121.340 77.540 ;
        RECT 121.970 77.370 125.050 77.540 ;
        RECT 125.680 77.370 128.760 77.540 ;
        RECT 129.390 77.370 132.470 77.540 ;
        RECT 133.100 77.370 136.180 77.540 ;
        RECT 22.150 76.300 37.000 76.500 ;
        RECT 22.150 74.350 22.350 76.300 ;
        RECT 22.760 75.620 23.800 75.790 ;
        RECT 26.355 75.620 36.395 75.790 ;
        RECT 23.970 75.060 24.140 75.560 ;
        RECT 26.015 75.060 26.185 75.560 ;
        RECT 22.760 74.830 23.800 75.000 ;
        RECT 26.355 74.830 36.395 75.000 ;
        RECT 36.800 74.350 37.000 76.300 ;
        RECT 22.150 74.150 37.000 74.350 ;
        RECT 22.200 73.050 36.950 73.250 ;
        RECT 22.200 69.700 22.400 73.050 ;
        RECT 22.710 72.490 23.750 72.660 ;
        RECT 26.400 72.490 36.440 72.660 ;
        RECT 23.965 71.930 24.135 72.430 ;
        RECT 26.015 71.930 26.185 72.430 ;
        RECT 22.710 71.700 23.750 71.870 ;
        RECT 26.400 71.700 36.440 71.870 ;
        RECT 23.965 71.140 24.135 71.640 ;
        RECT 26.015 71.140 26.185 71.640 ;
        RECT 22.710 70.910 23.750 71.080 ;
        RECT 26.400 70.910 36.440 71.080 ;
        RECT 23.965 70.350 24.135 70.850 ;
        RECT 26.015 70.350 26.185 70.850 ;
        RECT 22.710 70.120 23.750 70.290 ;
        RECT 26.400 70.120 36.440 70.290 ;
        RECT 36.750 69.700 36.950 73.050 ;
        RECT 22.200 69.500 36.950 69.700 ;
        RECT 40.450 71.150 104.350 71.550 ;
        RECT 40.450 57.050 40.850 71.150 ;
        RECT 48.280 70.510 50.820 70.680 ;
        RECT 51.420 70.510 57.710 70.680 ;
        RECT 58.310 70.510 64.600 70.680 ;
        RECT 65.200 70.510 71.490 70.680 ;
        RECT 72.090 70.510 78.380 70.680 ;
        RECT 78.980 70.510 85.270 70.680 ;
        RECT 85.870 70.510 88.410 70.680 ;
        RECT 47.895 69.450 48.065 70.450 ;
        RECT 51.035 69.450 51.205 70.450 ;
        RECT 57.925 69.450 58.095 70.450 ;
        RECT 64.815 69.450 64.985 70.450 ;
        RECT 71.705 69.450 71.875 70.450 ;
        RECT 78.595 69.450 78.765 70.450 ;
        RECT 85.485 69.450 85.655 70.450 ;
        RECT 88.625 69.450 88.795 70.450 ;
        RECT 48.280 69.220 50.820 69.390 ;
        RECT 51.420 69.220 57.710 69.390 ;
        RECT 58.310 69.220 64.600 69.390 ;
        RECT 65.200 69.220 71.490 69.390 ;
        RECT 72.090 69.220 78.380 69.390 ;
        RECT 78.980 69.220 85.270 69.390 ;
        RECT 85.870 69.220 88.410 69.390 ;
        RECT 47.895 68.160 48.065 69.160 ;
        RECT 51.035 68.160 51.205 69.160 ;
        RECT 57.925 68.160 58.095 69.160 ;
        RECT 64.815 68.160 64.985 69.160 ;
        RECT 71.705 68.160 71.875 69.160 ;
        RECT 78.595 68.160 78.765 69.160 ;
        RECT 85.485 68.160 85.655 69.160 ;
        RECT 88.625 68.160 88.795 69.160 ;
        RECT 48.280 67.930 50.820 68.100 ;
        RECT 51.420 67.930 57.710 68.100 ;
        RECT 58.310 67.930 64.600 68.100 ;
        RECT 65.200 67.930 71.490 68.100 ;
        RECT 72.090 67.930 78.380 68.100 ;
        RECT 78.980 67.930 85.270 68.100 ;
        RECT 85.870 67.930 88.410 68.100 ;
        RECT 47.895 66.870 48.065 67.870 ;
        RECT 51.035 66.870 51.205 67.870 ;
        RECT 57.925 66.870 58.095 67.870 ;
        RECT 64.815 66.870 64.985 67.870 ;
        RECT 71.705 66.870 71.875 67.870 ;
        RECT 78.595 66.870 78.765 67.870 ;
        RECT 85.485 66.870 85.655 67.870 ;
        RECT 88.625 66.870 88.795 67.870 ;
        RECT 48.280 66.640 50.820 66.810 ;
        RECT 51.420 66.640 57.710 66.810 ;
        RECT 58.310 66.640 64.600 66.810 ;
        RECT 65.200 66.640 71.490 66.810 ;
        RECT 72.090 66.640 78.380 66.810 ;
        RECT 78.980 66.640 85.270 66.810 ;
        RECT 85.870 66.640 88.410 66.810 ;
        RECT 47.895 65.580 48.065 66.580 ;
        RECT 51.035 65.580 51.205 66.580 ;
        RECT 57.925 65.580 58.095 66.580 ;
        RECT 64.815 65.580 64.985 66.580 ;
        RECT 71.705 65.580 71.875 66.580 ;
        RECT 78.595 65.580 78.765 66.580 ;
        RECT 85.485 65.580 85.655 66.580 ;
        RECT 88.625 65.580 88.795 66.580 ;
        RECT 95.850 66.250 96.250 71.150 ;
        RECT 98.320 70.440 101.360 70.610 ;
        RECT 97.935 69.880 98.105 70.380 ;
        RECT 98.320 69.650 101.360 69.820 ;
        RECT 99.280 68.980 102.320 69.150 ;
        RECT 98.895 68.420 99.065 68.920 ;
        RECT 99.280 68.190 102.320 68.360 ;
        RECT 103.950 66.250 104.350 71.150 ;
        RECT 95.850 65.850 104.350 66.250 ;
        RECT 48.280 65.350 50.820 65.520 ;
        RECT 51.420 65.350 57.710 65.520 ;
        RECT 58.310 65.350 64.600 65.520 ;
        RECT 65.200 65.350 71.490 65.520 ;
        RECT 72.090 65.350 78.380 65.520 ;
        RECT 78.980 65.350 85.270 65.520 ;
        RECT 85.870 65.350 88.410 65.520 ;
        RECT 47.895 64.290 48.065 65.290 ;
        RECT 51.035 64.290 51.205 65.290 ;
        RECT 57.925 64.290 58.095 65.290 ;
        RECT 64.815 64.290 64.985 65.290 ;
        RECT 71.705 64.290 71.875 65.290 ;
        RECT 78.595 64.290 78.765 65.290 ;
        RECT 85.485 64.290 85.655 65.290 ;
        RECT 88.625 64.290 88.795 65.290 ;
        RECT 48.280 64.060 50.820 64.230 ;
        RECT 51.420 64.060 57.710 64.230 ;
        RECT 58.310 64.060 64.600 64.230 ;
        RECT 65.200 64.060 71.490 64.230 ;
        RECT 72.090 64.060 78.380 64.230 ;
        RECT 78.980 64.060 85.270 64.230 ;
        RECT 85.870 64.060 88.410 64.230 ;
        RECT 47.895 63.000 48.065 64.000 ;
        RECT 51.035 63.000 51.205 64.000 ;
        RECT 57.925 63.000 58.095 64.000 ;
        RECT 64.815 63.000 64.985 64.000 ;
        RECT 71.705 63.000 71.875 64.000 ;
        RECT 78.595 63.000 78.765 64.000 ;
        RECT 85.485 63.000 85.655 64.000 ;
        RECT 88.625 63.000 88.795 64.000 ;
        RECT 48.280 62.770 50.820 62.940 ;
        RECT 51.420 62.770 57.710 62.940 ;
        RECT 58.310 62.770 64.600 62.940 ;
        RECT 65.200 62.770 71.490 62.940 ;
        RECT 72.090 62.770 78.380 62.940 ;
        RECT 78.980 62.770 85.270 62.940 ;
        RECT 85.870 62.770 88.410 62.940 ;
        RECT 47.895 61.710 48.065 62.710 ;
        RECT 51.035 61.710 51.205 62.710 ;
        RECT 57.925 61.710 58.095 62.710 ;
        RECT 64.815 61.710 64.985 62.710 ;
        RECT 71.705 61.710 71.875 62.710 ;
        RECT 78.595 61.710 78.765 62.710 ;
        RECT 85.485 61.710 85.655 62.710 ;
        RECT 88.625 61.710 88.795 62.710 ;
        RECT 48.280 61.480 50.820 61.650 ;
        RECT 51.420 61.480 57.710 61.650 ;
        RECT 58.310 61.480 64.600 61.650 ;
        RECT 65.200 61.480 71.490 61.650 ;
        RECT 72.090 61.480 78.380 61.650 ;
        RECT 78.980 61.480 85.270 61.650 ;
        RECT 85.870 61.480 88.410 61.650 ;
        RECT 47.895 60.420 48.065 61.420 ;
        RECT 51.035 60.420 51.205 61.420 ;
        RECT 57.925 60.420 58.095 61.420 ;
        RECT 64.815 60.420 64.985 61.420 ;
        RECT 71.705 60.420 71.875 61.420 ;
        RECT 78.595 60.420 78.765 61.420 ;
        RECT 85.485 60.420 85.655 61.420 ;
        RECT 88.625 60.420 88.795 61.420 ;
        RECT 48.280 60.190 50.820 60.360 ;
        RECT 51.420 60.190 57.710 60.360 ;
        RECT 58.310 60.190 64.600 60.360 ;
        RECT 65.200 60.190 71.490 60.360 ;
        RECT 72.090 60.190 78.380 60.360 ;
        RECT 78.980 60.190 85.270 60.360 ;
        RECT 85.870 60.190 88.410 60.360 ;
        RECT 95.850 57.050 96.250 65.850 ;
        RECT 40.450 56.650 96.250 57.050 ;
        RECT 40.450 42.700 40.850 56.650 ;
        RECT 41.580 56.030 66.620 56.200 ;
        RECT 70.080 56.030 95.120 56.200 ;
        RECT 41.195 54.970 41.365 55.970 ;
        RECT 66.835 54.970 67.005 55.970 ;
        RECT 69.695 54.970 69.865 55.970 ;
        RECT 95.335 54.970 95.505 55.970 ;
        RECT 41.580 54.740 66.620 54.910 ;
        RECT 70.080 54.740 95.120 54.910 ;
        RECT 41.195 53.680 41.365 54.680 ;
        RECT 66.835 53.680 67.005 54.680 ;
        RECT 69.695 53.680 69.865 54.680 ;
        RECT 95.335 53.680 95.505 54.680 ;
        RECT 41.580 53.450 66.620 53.620 ;
        RECT 70.080 53.450 95.120 53.620 ;
        RECT 41.195 52.390 41.365 53.390 ;
        RECT 66.835 52.390 67.005 53.390 ;
        RECT 69.695 52.390 69.865 53.390 ;
        RECT 95.335 52.390 95.505 53.390 ;
        RECT 41.580 52.160 66.620 52.330 ;
        RECT 70.080 52.160 95.120 52.330 ;
        RECT 41.195 51.100 41.365 52.100 ;
        RECT 66.835 51.100 67.005 52.100 ;
        RECT 69.695 51.100 69.865 52.100 ;
        RECT 95.335 51.100 95.505 52.100 ;
        RECT 41.580 50.870 66.620 51.040 ;
        RECT 70.080 50.870 95.120 51.040 ;
        RECT 41.195 49.810 41.365 50.810 ;
        RECT 66.835 49.810 67.005 50.810 ;
        RECT 69.695 49.810 69.865 50.810 ;
        RECT 95.335 49.810 95.505 50.810 ;
        RECT 41.580 49.580 66.620 49.750 ;
        RECT 70.080 49.580 95.120 49.750 ;
        RECT 41.195 48.520 41.365 49.520 ;
        RECT 66.835 48.520 67.005 49.520 ;
        RECT 69.695 48.520 69.865 49.520 ;
        RECT 95.335 48.520 95.505 49.520 ;
        RECT 41.580 48.290 66.620 48.460 ;
        RECT 70.080 48.290 95.120 48.460 ;
        RECT 41.195 47.230 41.365 48.230 ;
        RECT 66.835 47.230 67.005 48.230 ;
        RECT 69.695 47.230 69.865 48.230 ;
        RECT 95.335 47.230 95.505 48.230 ;
        RECT 41.580 47.000 66.620 47.170 ;
        RECT 70.080 47.000 95.120 47.170 ;
        RECT 41.195 45.940 41.365 46.940 ;
        RECT 66.835 45.940 67.005 46.940 ;
        RECT 69.695 45.940 69.865 46.940 ;
        RECT 95.335 45.940 95.505 46.940 ;
        RECT 41.580 45.710 66.620 45.880 ;
        RECT 70.080 45.710 95.120 45.880 ;
        RECT 41.195 44.650 41.365 45.650 ;
        RECT 66.835 44.650 67.005 45.650 ;
        RECT 69.695 44.650 69.865 45.650 ;
        RECT 95.335 44.650 95.505 45.650 ;
        RECT 41.580 44.420 66.620 44.590 ;
        RECT 70.080 44.420 95.120 44.590 ;
        RECT 41.195 43.360 41.365 44.360 ;
        RECT 66.835 43.360 67.005 44.360 ;
        RECT 69.695 43.360 69.865 44.360 ;
        RECT 95.335 43.360 95.505 44.360 ;
        RECT 41.580 43.130 66.620 43.300 ;
        RECT 70.080 43.130 95.120 43.300 ;
        RECT 95.850 42.700 96.250 56.650 ;
        RECT 40.450 42.300 96.250 42.700 ;
        RECT 97.250 64.450 104.700 64.850 ;
        RECT 97.250 41.300 97.650 64.450 ;
        RECT 98.370 63.500 99.410 63.670 ;
        RECT 100.270 63.500 101.310 63.670 ;
        RECT 98.030 62.940 98.200 63.440 ;
        RECT 99.930 62.940 100.100 63.440 ;
        RECT 98.370 62.710 99.410 62.880 ;
        RECT 100.270 62.710 101.310 62.880 ;
        RECT 98.540 60.580 99.540 60.750 ;
        RECT 99.830 60.580 100.830 60.750 ;
        RECT 101.120 60.580 102.120 60.750 ;
        RECT 102.410 60.580 103.410 60.750 ;
        RECT 98.310 42.870 98.480 60.410 ;
        RECT 99.600 42.870 99.770 60.410 ;
        RECT 100.890 42.870 101.060 60.410 ;
        RECT 102.180 42.870 102.350 60.410 ;
        RECT 103.470 42.870 103.640 60.410 ;
        RECT 98.540 42.530 99.540 42.700 ;
        RECT 99.830 42.530 100.830 42.700 ;
        RECT 101.120 42.530 102.120 42.700 ;
        RECT 102.410 42.530 103.410 42.700 ;
        RECT 40.450 40.900 97.650 41.300 ;
        RECT 40.450 36.900 40.850 40.900 ;
        RECT 44.455 40.090 48.995 40.260 ;
        RECT 49.505 40.090 58.545 40.260 ;
        RECT 59.055 40.090 68.095 40.260 ;
        RECT 68.605 40.090 77.645 40.260 ;
        RECT 78.155 40.090 87.195 40.260 ;
        RECT 87.705 40.090 92.245 40.260 ;
        RECT 44.115 39.030 44.285 40.030 ;
        RECT 49.165 39.030 49.335 40.030 ;
        RECT 58.715 39.030 58.885 40.030 ;
        RECT 68.265 39.030 68.435 40.030 ;
        RECT 77.815 39.030 77.985 40.030 ;
        RECT 87.365 39.030 87.535 40.030 ;
        RECT 92.415 39.030 92.585 40.030 ;
        RECT 44.455 38.800 48.995 38.970 ;
        RECT 49.505 38.800 58.545 38.970 ;
        RECT 59.055 38.800 68.095 38.970 ;
        RECT 68.605 38.800 77.645 38.970 ;
        RECT 78.155 38.800 87.195 38.970 ;
        RECT 87.705 38.800 92.245 38.970 ;
        RECT 44.115 37.740 44.285 38.740 ;
        RECT 49.165 37.740 49.335 38.740 ;
        RECT 58.715 37.740 58.885 38.740 ;
        RECT 68.265 37.740 68.435 38.740 ;
        RECT 77.815 37.740 77.985 38.740 ;
        RECT 87.365 37.740 87.535 38.740 ;
        RECT 92.415 37.740 92.585 38.740 ;
        RECT 44.455 37.510 48.995 37.680 ;
        RECT 49.505 37.510 58.545 37.680 ;
        RECT 59.055 37.510 68.095 37.680 ;
        RECT 68.605 37.510 77.645 37.680 ;
        RECT 78.155 37.510 87.195 37.680 ;
        RECT 87.705 37.510 92.245 37.680 ;
        RECT 104.300 36.900 104.700 64.450 ;
        RECT 107.410 60.770 107.580 76.810 ;
        RECT 108.200 60.770 108.370 76.810 ;
        RECT 108.990 60.770 109.160 76.810 ;
        RECT 109.780 60.770 109.950 76.810 ;
        RECT 111.110 60.780 111.280 76.820 ;
        RECT 111.900 60.780 112.070 76.820 ;
        RECT 112.690 60.780 112.860 76.820 ;
        RECT 113.480 60.780 113.650 76.820 ;
        RECT 114.820 60.780 114.990 76.820 ;
        RECT 115.610 60.780 115.780 76.820 ;
        RECT 116.400 60.780 116.570 76.820 ;
        RECT 117.190 60.780 117.360 76.820 ;
        RECT 118.530 60.780 118.700 76.820 ;
        RECT 119.320 60.780 119.490 76.820 ;
        RECT 120.110 60.780 120.280 76.820 ;
        RECT 120.900 60.780 121.070 76.820 ;
        RECT 122.240 60.780 122.410 76.820 ;
        RECT 123.030 60.780 123.200 76.820 ;
        RECT 123.820 60.780 123.990 76.820 ;
        RECT 124.610 60.780 124.780 76.820 ;
        RECT 125.950 60.780 126.120 76.820 ;
        RECT 126.740 60.780 126.910 76.820 ;
        RECT 127.530 60.780 127.700 76.820 ;
        RECT 128.320 60.780 128.490 76.820 ;
        RECT 129.660 60.780 129.830 76.820 ;
        RECT 130.450 60.780 130.620 76.820 ;
        RECT 131.240 60.780 131.410 76.820 ;
        RECT 132.030 60.780 132.200 76.820 ;
        RECT 133.370 60.780 133.540 76.820 ;
        RECT 134.160 60.780 134.330 76.820 ;
        RECT 134.950 60.780 135.120 76.820 ;
        RECT 135.740 60.780 135.910 76.820 ;
        RECT 107.640 60.385 108.140 60.555 ;
        RECT 108.430 60.385 108.930 60.555 ;
        RECT 109.220 60.385 109.720 60.555 ;
        RECT 111.340 60.395 111.840 60.565 ;
        RECT 112.130 60.395 112.630 60.565 ;
        RECT 112.920 60.395 113.420 60.565 ;
        RECT 115.050 60.395 115.550 60.565 ;
        RECT 115.840 60.395 116.340 60.565 ;
        RECT 116.630 60.395 117.130 60.565 ;
        RECT 118.760 60.395 119.260 60.565 ;
        RECT 119.550 60.395 120.050 60.565 ;
        RECT 120.340 60.395 120.840 60.565 ;
        RECT 122.470 60.395 122.970 60.565 ;
        RECT 123.260 60.395 123.760 60.565 ;
        RECT 124.050 60.395 124.550 60.565 ;
        RECT 126.180 60.395 126.680 60.565 ;
        RECT 126.970 60.395 127.470 60.565 ;
        RECT 127.760 60.395 128.260 60.565 ;
        RECT 129.890 60.395 130.390 60.565 ;
        RECT 130.680 60.395 131.180 60.565 ;
        RECT 131.470 60.395 131.970 60.565 ;
        RECT 133.600 60.395 134.100 60.565 ;
        RECT 134.390 60.395 134.890 60.565 ;
        RECT 135.180 60.395 135.680 60.565 ;
        RECT 107.140 59.690 110.220 59.860 ;
        RECT 110.840 59.700 113.920 59.870 ;
        RECT 114.550 59.700 117.630 59.870 ;
        RECT 118.260 59.700 121.340 59.870 ;
        RECT 121.970 59.700 125.050 59.870 ;
        RECT 125.680 59.700 128.760 59.870 ;
        RECT 129.390 59.700 132.470 59.870 ;
        RECT 133.100 59.700 136.180 59.870 ;
        RECT 107.140 58.310 110.220 58.480 ;
        RECT 110.840 58.320 113.920 58.490 ;
        RECT 114.550 58.320 117.630 58.490 ;
        RECT 118.260 58.320 121.340 58.490 ;
        RECT 121.970 58.320 125.050 58.490 ;
        RECT 125.680 58.320 128.760 58.490 ;
        RECT 129.390 58.320 132.470 58.490 ;
        RECT 133.100 58.320 136.180 58.490 ;
        RECT 107.640 57.620 109.720 57.790 ;
        RECT 111.340 57.630 113.420 57.800 ;
        RECT 115.050 57.630 117.130 57.800 ;
        RECT 118.760 57.630 120.840 57.800 ;
        RECT 122.470 57.630 124.550 57.800 ;
        RECT 126.180 57.630 128.260 57.800 ;
        RECT 129.890 57.630 131.970 57.800 ;
        RECT 133.600 57.630 135.680 57.800 ;
        RECT 107.410 50.410 107.580 57.450 ;
        RECT 108.200 50.410 108.370 57.450 ;
        RECT 108.990 50.410 109.160 57.450 ;
        RECT 109.780 50.410 109.950 57.450 ;
        RECT 111.110 50.420 111.280 57.460 ;
        RECT 111.900 50.420 112.070 57.460 ;
        RECT 112.690 50.420 112.860 57.460 ;
        RECT 113.480 50.420 113.650 57.460 ;
        RECT 114.820 50.420 114.990 57.460 ;
        RECT 115.610 50.420 115.780 57.460 ;
        RECT 116.400 50.420 116.570 57.460 ;
        RECT 117.190 50.420 117.360 57.460 ;
        RECT 118.530 50.420 118.700 57.460 ;
        RECT 119.320 50.420 119.490 57.460 ;
        RECT 120.110 50.420 120.280 57.460 ;
        RECT 120.900 50.420 121.070 57.460 ;
        RECT 122.240 50.420 122.410 57.460 ;
        RECT 123.030 50.420 123.200 57.460 ;
        RECT 123.820 50.420 123.990 57.460 ;
        RECT 124.610 50.420 124.780 57.460 ;
        RECT 125.950 50.420 126.120 57.460 ;
        RECT 126.740 50.420 126.910 57.460 ;
        RECT 127.530 50.420 127.700 57.460 ;
        RECT 128.320 50.420 128.490 57.460 ;
        RECT 129.660 50.420 129.830 57.460 ;
        RECT 130.450 50.420 130.620 57.460 ;
        RECT 131.240 50.420 131.410 57.460 ;
        RECT 132.030 50.420 132.200 57.460 ;
        RECT 133.370 50.420 133.540 57.460 ;
        RECT 134.160 50.420 134.330 57.460 ;
        RECT 134.950 50.420 135.120 57.460 ;
        RECT 135.740 50.420 135.910 57.460 ;
        RECT 107.140 49.690 110.220 49.860 ;
        RECT 110.840 49.700 113.920 49.870 ;
        RECT 114.550 49.700 117.630 49.870 ;
        RECT 118.260 49.700 121.340 49.870 ;
        RECT 121.970 49.700 125.050 49.870 ;
        RECT 125.680 49.700 128.760 49.870 ;
        RECT 129.390 49.700 132.470 49.870 ;
        RECT 133.100 49.700 136.180 49.870 ;
        RECT 40.450 36.500 104.700 36.900 ;
        RECT 105.200 35.580 105.370 47.240 ;
        RECT 105.850 44.830 106.540 46.990 ;
        RECT 107.020 44.830 107.710 46.990 ;
        RECT 108.190 44.830 108.880 46.990 ;
        RECT 109.360 44.830 110.050 46.990 ;
        RECT 110.530 44.830 111.220 46.990 ;
        RECT 111.700 44.830 112.390 46.990 ;
        RECT 112.870 44.830 113.560 46.990 ;
        RECT 114.040 44.830 114.730 46.990 ;
        RECT 115.210 44.830 115.900 46.990 ;
        RECT 116.380 44.830 117.070 46.990 ;
        RECT 117.550 44.830 118.240 46.990 ;
        RECT 118.720 44.830 119.410 46.990 ;
        RECT 119.890 44.830 120.580 46.990 ;
        RECT 121.060 44.830 121.750 46.990 ;
        RECT 122.230 44.830 122.920 46.990 ;
        RECT 123.400 44.830 124.090 46.990 ;
        RECT 124.570 44.830 125.260 46.990 ;
        RECT 125.740 44.830 126.430 46.990 ;
        RECT 126.910 44.830 127.600 46.990 ;
        RECT 128.080 44.830 128.770 46.990 ;
        RECT 129.250 44.830 129.940 46.990 ;
        RECT 130.420 44.830 131.110 46.990 ;
        RECT 131.590 44.830 132.280 46.990 ;
        RECT 132.760 44.830 133.450 46.990 ;
        RECT 133.930 44.830 134.620 46.990 ;
        RECT 135.100 44.830 135.790 46.990 ;
        RECT 136.270 44.830 136.960 46.990 ;
        RECT 105.850 35.830 106.540 37.990 ;
        RECT 107.020 35.830 107.710 37.990 ;
        RECT 108.190 35.830 108.880 37.990 ;
        RECT 109.360 35.830 110.050 37.990 ;
        RECT 110.530 35.830 111.220 37.990 ;
        RECT 111.700 35.830 112.390 37.990 ;
        RECT 112.870 35.830 113.560 37.990 ;
        RECT 114.040 35.830 114.730 37.990 ;
        RECT 115.210 35.830 115.900 37.990 ;
        RECT 116.380 35.830 117.070 37.990 ;
        RECT 117.550 35.830 118.240 37.990 ;
        RECT 118.720 35.830 119.410 37.990 ;
        RECT 119.890 35.830 120.580 37.990 ;
        RECT 121.060 35.830 121.750 37.990 ;
        RECT 122.230 35.830 122.920 37.990 ;
        RECT 123.400 35.830 124.090 37.990 ;
        RECT 124.570 35.830 125.260 37.990 ;
        RECT 125.740 35.830 126.430 37.990 ;
        RECT 126.910 35.830 127.600 37.990 ;
        RECT 128.080 35.830 128.770 37.990 ;
        RECT 129.250 35.830 129.940 37.990 ;
        RECT 130.420 35.830 131.110 37.990 ;
        RECT 131.590 35.830 132.280 37.990 ;
        RECT 132.760 35.830 133.450 37.990 ;
        RECT 133.930 35.830 134.620 37.990 ;
        RECT 135.100 35.830 135.790 37.990 ;
        RECT 136.270 35.830 136.960 37.990 ;
        RECT 137.440 35.580 137.610 47.240 ;
        RECT 105.600 35.180 137.210 35.350 ;
        RECT 20.500 31.000 95.100 31.400 ;
        RECT 20.500 23.300 20.900 31.000 ;
        RECT 21.630 30.370 22.670 30.540 ;
        RECT 23.270 30.370 32.310 30.540 ;
        RECT 32.910 30.370 41.950 30.540 ;
        RECT 42.550 30.370 51.590 30.540 ;
        RECT 52.190 30.370 61.230 30.540 ;
        RECT 61.830 30.370 70.870 30.540 ;
        RECT 71.470 30.370 80.510 30.540 ;
        RECT 81.110 30.370 82.150 30.540 ;
        RECT 21.245 27.310 21.415 30.310 ;
        RECT 22.885 27.310 23.055 30.310 ;
        RECT 32.525 27.310 32.695 30.310 ;
        RECT 42.165 27.310 42.335 30.310 ;
        RECT 51.805 27.310 51.975 30.310 ;
        RECT 61.445 27.310 61.615 30.310 ;
        RECT 71.085 27.310 71.255 30.310 ;
        RECT 80.725 27.310 80.895 30.310 ;
        RECT 82.365 27.310 82.535 30.310 ;
        RECT 82.900 28.400 83.300 31.000 ;
        RECT 84.020 30.385 94.020 30.555 ;
        RECT 83.790 29.130 83.960 30.170 ;
        RECT 94.080 29.130 94.250 30.170 ;
        RECT 84.020 28.745 94.020 28.915 ;
        RECT 94.700 28.400 95.100 31.000 ;
        RECT 82.900 28.000 95.100 28.400 ;
        RECT 96.250 31.000 133.100 31.400 ;
        RECT 21.630 27.080 22.670 27.250 ;
        RECT 23.270 27.080 32.310 27.250 ;
        RECT 32.910 27.080 41.950 27.250 ;
        RECT 42.550 27.080 51.590 27.250 ;
        RECT 52.190 27.080 61.230 27.250 ;
        RECT 61.830 27.080 70.870 27.250 ;
        RECT 71.470 27.080 80.510 27.250 ;
        RECT 81.110 27.080 82.150 27.250 ;
        RECT 21.245 24.020 21.415 27.020 ;
        RECT 22.885 24.020 23.055 27.020 ;
        RECT 32.525 24.020 32.695 27.020 ;
        RECT 42.165 24.020 42.335 27.020 ;
        RECT 51.805 24.020 51.975 27.020 ;
        RECT 61.445 24.020 61.615 27.020 ;
        RECT 71.085 24.020 71.255 27.020 ;
        RECT 80.725 24.020 80.895 27.020 ;
        RECT 82.365 24.020 82.535 27.020 ;
        RECT 21.630 23.790 22.670 23.960 ;
        RECT 23.270 23.790 32.310 23.960 ;
        RECT 32.910 23.790 41.950 23.960 ;
        RECT 42.550 23.790 51.590 23.960 ;
        RECT 52.190 23.790 61.230 23.960 ;
        RECT 61.830 23.790 70.870 23.960 ;
        RECT 71.470 23.790 80.510 23.960 ;
        RECT 81.110 23.790 82.150 23.960 ;
        RECT 82.900 23.300 83.300 28.000 ;
        RECT 96.250 26.900 96.650 31.000 ;
        RECT 97.490 30.380 98.490 30.550 ;
        RECT 99.920 30.290 100.960 30.460 ;
        RECT 101.470 30.290 104.510 30.460 ;
        RECT 105.020 30.290 108.060 30.460 ;
        RECT 108.570 30.290 111.610 30.460 ;
        RECT 112.120 30.290 115.160 30.460 ;
        RECT 115.670 30.290 116.710 30.460 ;
        RECT 20.500 22.900 83.300 23.300 ;
        RECT 84.300 26.500 96.650 26.900 ;
        RECT 84.300 22.650 84.700 26.500 ;
        RECT 85.470 25.790 95.510 25.960 ;
        RECT 85.130 24.730 85.300 25.730 ;
        RECT 95.680 24.730 95.850 25.730 ;
        RECT 97.260 25.170 97.430 30.210 ;
        RECT 98.550 25.170 98.720 30.210 ;
        RECT 99.580 27.230 99.750 30.230 ;
        RECT 101.130 27.230 101.300 30.230 ;
        RECT 104.680 27.230 104.850 30.230 ;
        RECT 108.230 27.230 108.400 30.230 ;
        RECT 111.780 27.230 111.950 30.230 ;
        RECT 115.330 27.230 115.500 30.230 ;
        RECT 116.880 27.230 117.050 30.230 ;
        RECT 117.650 28.970 119.810 30.380 ;
        RECT 129.950 28.970 132.110 30.380 ;
        RECT 99.920 27.000 100.960 27.170 ;
        RECT 101.470 27.000 104.510 27.170 ;
        RECT 105.020 27.000 108.060 27.170 ;
        RECT 108.570 27.000 111.610 27.170 ;
        RECT 112.120 27.000 115.160 27.170 ;
        RECT 115.670 27.000 116.710 27.170 ;
        RECT 117.650 27.080 119.810 28.490 ;
        RECT 129.950 27.080 132.110 28.490 ;
        RECT 97.490 24.830 98.490 25.000 ;
        RECT 85.470 24.500 95.510 24.670 ;
        RECT 85.130 23.440 85.300 24.440 ;
        RECT 95.680 23.440 95.850 24.440 ;
        RECT 99.580 23.940 99.750 26.940 ;
        RECT 101.130 23.940 101.300 26.940 ;
        RECT 104.680 23.940 104.850 26.940 ;
        RECT 108.230 23.940 108.400 26.940 ;
        RECT 111.780 23.940 111.950 26.940 ;
        RECT 115.330 23.940 115.500 26.940 ;
        RECT 116.880 23.940 117.050 26.940 ;
        RECT 117.650 25.190 119.810 26.600 ;
        RECT 129.950 25.190 132.110 26.600 ;
        RECT 99.920 23.710 100.960 23.880 ;
        RECT 101.470 23.710 104.510 23.880 ;
        RECT 105.020 23.710 108.060 23.880 ;
        RECT 108.570 23.710 111.610 23.880 ;
        RECT 112.120 23.710 115.160 23.880 ;
        RECT 115.670 23.710 116.710 23.880 ;
        RECT 85.470 23.210 95.510 23.380 ;
        RECT 117.650 23.300 119.810 24.710 ;
        RECT 129.950 23.300 132.110 24.710 ;
        RECT 132.700 22.650 133.100 31.000 ;
        RECT 84.300 22.250 133.100 22.650 ;
        RECT 20.500 17.150 134.150 17.550 ;
        RECT 20.500 5.500 20.900 17.150 ;
        RECT 21.630 16.380 22.670 16.550 ;
        RECT 23.180 16.380 38.220 16.550 ;
        RECT 38.730 16.380 53.770 16.550 ;
        RECT 54.280 16.380 69.320 16.550 ;
        RECT 69.830 16.380 84.870 16.550 ;
        RECT 85.380 16.380 100.420 16.550 ;
        RECT 100.930 16.380 115.970 16.550 ;
        RECT 116.480 16.380 131.520 16.550 ;
        RECT 132.030 16.380 133.070 16.550 ;
        RECT 21.290 15.320 21.460 16.320 ;
        RECT 22.840 15.320 23.010 16.320 ;
        RECT 38.390 15.320 38.560 16.320 ;
        RECT 53.940 15.320 54.110 16.320 ;
        RECT 69.490 15.320 69.660 16.320 ;
        RECT 85.040 15.320 85.210 16.320 ;
        RECT 100.590 15.320 100.760 16.320 ;
        RECT 116.140 15.320 116.310 16.320 ;
        RECT 131.690 15.320 131.860 16.320 ;
        RECT 133.240 15.320 133.410 16.320 ;
        RECT 21.630 15.090 22.670 15.260 ;
        RECT 23.180 15.090 38.220 15.260 ;
        RECT 38.730 15.090 53.770 15.260 ;
        RECT 54.280 15.090 69.320 15.260 ;
        RECT 69.830 15.090 84.870 15.260 ;
        RECT 85.380 15.090 100.420 15.260 ;
        RECT 100.930 15.090 115.970 15.260 ;
        RECT 116.480 15.090 131.520 15.260 ;
        RECT 132.030 15.090 133.070 15.260 ;
        RECT 21.290 14.030 21.460 15.030 ;
        RECT 22.840 14.030 23.010 15.030 ;
        RECT 38.390 14.030 38.560 15.030 ;
        RECT 53.940 14.030 54.110 15.030 ;
        RECT 69.490 14.030 69.660 15.030 ;
        RECT 85.040 14.030 85.210 15.030 ;
        RECT 100.590 14.030 100.760 15.030 ;
        RECT 116.140 14.030 116.310 15.030 ;
        RECT 131.690 14.030 131.860 15.030 ;
        RECT 133.240 14.030 133.410 15.030 ;
        RECT 21.630 13.800 22.670 13.970 ;
        RECT 23.180 13.800 38.220 13.970 ;
        RECT 38.730 13.800 53.770 13.970 ;
        RECT 54.280 13.800 69.320 13.970 ;
        RECT 69.830 13.800 84.870 13.970 ;
        RECT 85.380 13.800 100.420 13.970 ;
        RECT 100.930 13.800 115.970 13.970 ;
        RECT 116.480 13.800 131.520 13.970 ;
        RECT 132.030 13.800 133.070 13.970 ;
        RECT 21.290 12.740 21.460 13.740 ;
        RECT 22.840 12.740 23.010 13.740 ;
        RECT 38.390 12.740 38.560 13.740 ;
        RECT 53.940 12.740 54.110 13.740 ;
        RECT 69.490 12.740 69.660 13.740 ;
        RECT 85.040 12.740 85.210 13.740 ;
        RECT 100.590 12.740 100.760 13.740 ;
        RECT 116.140 12.740 116.310 13.740 ;
        RECT 131.690 12.740 131.860 13.740 ;
        RECT 133.240 12.740 133.410 13.740 ;
        RECT 21.630 12.510 22.670 12.680 ;
        RECT 23.180 12.510 38.220 12.680 ;
        RECT 38.730 12.510 53.770 12.680 ;
        RECT 54.280 12.510 69.320 12.680 ;
        RECT 69.830 12.510 84.870 12.680 ;
        RECT 85.380 12.510 100.420 12.680 ;
        RECT 100.930 12.510 115.970 12.680 ;
        RECT 116.480 12.510 131.520 12.680 ;
        RECT 132.030 12.510 133.070 12.680 ;
        RECT 21.290 11.450 21.460 12.450 ;
        RECT 22.840 11.450 23.010 12.450 ;
        RECT 38.390 11.450 38.560 12.450 ;
        RECT 53.940 11.450 54.110 12.450 ;
        RECT 69.490 11.450 69.660 12.450 ;
        RECT 85.040 11.450 85.210 12.450 ;
        RECT 100.590 11.450 100.760 12.450 ;
        RECT 116.140 11.450 116.310 12.450 ;
        RECT 131.690 11.450 131.860 12.450 ;
        RECT 133.240 11.450 133.410 12.450 ;
        RECT 21.630 11.220 22.670 11.390 ;
        RECT 23.180 11.220 38.220 11.390 ;
        RECT 38.730 11.220 53.770 11.390 ;
        RECT 54.280 11.220 69.320 11.390 ;
        RECT 69.830 11.220 84.870 11.390 ;
        RECT 85.380 11.220 100.420 11.390 ;
        RECT 100.930 11.220 115.970 11.390 ;
        RECT 116.480 11.220 131.520 11.390 ;
        RECT 132.030 11.220 133.070 11.390 ;
        RECT 21.290 10.160 21.460 11.160 ;
        RECT 22.840 10.160 23.010 11.160 ;
        RECT 38.390 10.160 38.560 11.160 ;
        RECT 53.940 10.160 54.110 11.160 ;
        RECT 69.490 10.160 69.660 11.160 ;
        RECT 85.040 10.160 85.210 11.160 ;
        RECT 100.590 10.160 100.760 11.160 ;
        RECT 116.140 10.160 116.310 11.160 ;
        RECT 131.690 10.160 131.860 11.160 ;
        RECT 133.240 10.160 133.410 11.160 ;
        RECT 21.630 9.930 22.670 10.100 ;
        RECT 23.180 9.930 38.220 10.100 ;
        RECT 38.730 9.930 53.770 10.100 ;
        RECT 54.280 9.930 69.320 10.100 ;
        RECT 69.830 9.930 84.870 10.100 ;
        RECT 85.380 9.930 100.420 10.100 ;
        RECT 100.930 9.930 115.970 10.100 ;
        RECT 116.480 9.930 131.520 10.100 ;
        RECT 132.030 9.930 133.070 10.100 ;
        RECT 21.290 8.870 21.460 9.870 ;
        RECT 22.840 8.870 23.010 9.870 ;
        RECT 38.390 8.870 38.560 9.870 ;
        RECT 53.940 8.870 54.110 9.870 ;
        RECT 69.490 8.870 69.660 9.870 ;
        RECT 85.040 8.870 85.210 9.870 ;
        RECT 100.590 8.870 100.760 9.870 ;
        RECT 116.140 8.870 116.310 9.870 ;
        RECT 131.690 8.870 131.860 9.870 ;
        RECT 133.240 8.870 133.410 9.870 ;
        RECT 21.630 8.640 22.670 8.810 ;
        RECT 23.180 8.640 38.220 8.810 ;
        RECT 38.730 8.640 53.770 8.810 ;
        RECT 54.280 8.640 69.320 8.810 ;
        RECT 69.830 8.640 84.870 8.810 ;
        RECT 85.380 8.640 100.420 8.810 ;
        RECT 100.930 8.640 115.970 8.810 ;
        RECT 116.480 8.640 131.520 8.810 ;
        RECT 132.030 8.640 133.070 8.810 ;
        RECT 21.290 7.580 21.460 8.580 ;
        RECT 22.840 7.580 23.010 8.580 ;
        RECT 38.390 7.580 38.560 8.580 ;
        RECT 53.940 7.580 54.110 8.580 ;
        RECT 69.490 7.580 69.660 8.580 ;
        RECT 85.040 7.580 85.210 8.580 ;
        RECT 100.590 7.580 100.760 8.580 ;
        RECT 116.140 7.580 116.310 8.580 ;
        RECT 131.690 7.580 131.860 8.580 ;
        RECT 133.240 7.580 133.410 8.580 ;
        RECT 21.630 7.350 22.670 7.520 ;
        RECT 23.180 7.350 38.220 7.520 ;
        RECT 38.730 7.350 53.770 7.520 ;
        RECT 54.280 7.350 69.320 7.520 ;
        RECT 69.830 7.350 84.870 7.520 ;
        RECT 85.380 7.350 100.420 7.520 ;
        RECT 100.930 7.350 115.970 7.520 ;
        RECT 116.480 7.350 131.520 7.520 ;
        RECT 132.030 7.350 133.070 7.520 ;
        RECT 21.290 6.290 21.460 7.290 ;
        RECT 22.840 6.290 23.010 7.290 ;
        RECT 38.390 6.290 38.560 7.290 ;
        RECT 53.940 6.290 54.110 7.290 ;
        RECT 69.490 6.290 69.660 7.290 ;
        RECT 85.040 6.290 85.210 7.290 ;
        RECT 100.590 6.290 100.760 7.290 ;
        RECT 116.140 6.290 116.310 7.290 ;
        RECT 131.690 6.290 131.860 7.290 ;
        RECT 133.240 6.290 133.410 7.290 ;
        RECT 21.630 6.060 22.670 6.230 ;
        RECT 23.180 6.060 38.220 6.230 ;
        RECT 38.730 6.060 53.770 6.230 ;
        RECT 54.280 6.060 69.320 6.230 ;
        RECT 69.830 6.060 84.870 6.230 ;
        RECT 85.380 6.060 100.420 6.230 ;
        RECT 100.930 6.060 115.970 6.230 ;
        RECT 116.480 6.060 131.520 6.230 ;
        RECT 132.030 6.060 133.070 6.230 ;
        RECT 133.750 5.500 134.150 17.150 ;
        RECT 20.500 5.100 134.150 5.500 ;
      LAYER met1 ;
        RECT 35.190 155.920 109.250 156.400 ;
        RECT 75.295 155.720 75.585 155.765 ;
        RECT 76.200 155.720 76.520 155.780 ;
        RECT 75.295 155.580 76.520 155.720 ;
        RECT 75.295 155.535 75.585 155.580 ;
        RECT 76.200 155.520 76.520 155.580 ;
        RECT 37.560 154.500 37.880 154.760 ;
        RECT 74.820 154.500 75.140 154.760 ;
        RECT 38.495 154.020 38.785 154.065 ;
        RECT 51.820 154.020 52.140 154.080 ;
        RECT 55.500 154.020 55.820 154.080 ;
        RECT 38.495 153.880 55.820 154.020 ;
        RECT 38.495 153.835 38.785 153.880 ;
        RECT 51.820 153.820 52.140 153.880 ;
        RECT 55.500 153.820 55.820 153.880 ;
        RECT 35.190 153.200 110.030 153.680 ;
        RECT 54.580 153.000 54.900 153.060 ;
        RECT 58.735 153.000 59.025 153.045 ;
        RECT 54.580 152.860 59.025 153.000 ;
        RECT 54.580 152.800 54.900 152.860 ;
        RECT 58.735 152.815 59.025 152.860 ;
        RECT 60.560 153.000 60.880 153.060 ;
        RECT 63.335 153.000 63.625 153.045 ;
        RECT 60.560 152.860 63.625 153.000 ;
        RECT 60.560 152.800 60.880 152.860 ;
        RECT 63.335 152.815 63.625 152.860 ;
        RECT 65.175 153.000 65.465 153.045 ;
        RECT 68.380 153.000 68.700 153.060 ;
        RECT 65.175 152.860 68.700 153.000 ;
        RECT 65.175 152.815 65.465 152.860 ;
        RECT 68.380 152.800 68.700 152.860 ;
        RECT 76.290 152.860 87.470 153.000 ;
        RECT 56.895 152.660 57.185 152.705 ;
        RECT 67.920 152.660 68.240 152.720 ;
        RECT 56.895 152.520 68.240 152.660 ;
        RECT 56.895 152.475 57.185 152.520 ;
        RECT 55.500 152.120 55.820 152.380 ;
        RECT 59.195 152.320 59.485 152.365 ;
        RECT 61.480 152.320 61.800 152.380 ;
        RECT 62.490 152.365 62.630 152.520 ;
        RECT 67.920 152.460 68.240 152.520 ;
        RECT 69.755 152.660 70.405 152.705 ;
        RECT 71.140 152.660 71.460 152.720 ;
        RECT 73.355 152.660 73.645 152.705 ;
        RECT 69.755 152.520 73.645 152.660 ;
        RECT 69.755 152.475 70.405 152.520 ;
        RECT 71.140 152.460 71.460 152.520 ;
        RECT 73.055 152.475 73.645 152.520 ;
        RECT 59.195 152.180 61.800 152.320 ;
        RECT 59.195 152.135 59.485 152.180 ;
        RECT 61.480 152.120 61.800 152.180 ;
        RECT 62.415 152.135 62.705 152.365 ;
        RECT 63.780 152.120 64.100 152.380 ;
        RECT 64.240 152.320 64.560 152.380 ;
        RECT 64.715 152.320 65.005 152.365 ;
        RECT 64.240 152.180 65.005 152.320 ;
        RECT 64.240 152.120 64.560 152.180 ;
        RECT 64.715 152.135 65.005 152.180 ;
        RECT 66.560 152.320 66.850 152.365 ;
        RECT 68.395 152.320 68.685 152.365 ;
        RECT 71.975 152.320 72.265 152.365 ;
        RECT 66.560 152.180 72.265 152.320 ;
        RECT 66.560 152.135 66.850 152.180 ;
        RECT 68.395 152.135 68.685 152.180 ;
        RECT 71.975 152.135 72.265 152.180 ;
        RECT 73.055 152.160 73.345 152.475 ;
        RECT 76.290 152.365 76.430 152.860 ;
        RECT 79.875 152.660 80.525 152.705 ;
        RECT 83.475 152.660 83.765 152.705 ;
        RECT 85.875 152.660 86.165 152.705 ;
        RECT 79.875 152.520 86.165 152.660 ;
        RECT 79.875 152.475 80.525 152.520 ;
        RECT 83.175 152.475 83.765 152.520 ;
        RECT 85.875 152.475 86.165 152.520 ;
        RECT 76.215 152.135 76.505 152.365 ;
        RECT 76.680 152.320 76.970 152.365 ;
        RECT 78.515 152.320 78.805 152.365 ;
        RECT 82.095 152.320 82.385 152.365 ;
        RECT 76.680 152.180 82.385 152.320 ;
        RECT 76.680 152.135 76.970 152.180 ;
        RECT 78.515 152.135 78.805 152.180 ;
        RECT 82.095 152.135 82.385 152.180 ;
        RECT 83.175 152.160 83.465 152.475 ;
        RECT 87.330 152.380 87.470 152.860 ;
        RECT 91.380 152.705 91.700 152.720 ;
        RECT 90.915 152.660 91.700 152.705 ;
        RECT 94.515 152.660 94.805 152.705 ;
        RECT 90.915 152.520 94.805 152.660 ;
        RECT 90.915 152.475 91.700 152.520 ;
        RECT 91.380 152.460 91.700 152.475 ;
        RECT 94.215 152.475 94.805 152.520 ;
        RECT 86.320 152.320 86.640 152.380 ;
        RECT 83.650 152.180 86.640 152.320 ;
        RECT 56.880 151.980 57.200 152.040 ;
        RECT 66.095 151.980 66.385 152.025 ;
        RECT 56.880 151.840 66.385 151.980 ;
        RECT 56.880 151.780 57.200 151.840 ;
        RECT 66.095 151.795 66.385 151.840 ;
        RECT 67.460 151.780 67.780 152.040 ;
        RECT 77.580 151.780 77.900 152.040 ;
        RECT 66.965 151.640 67.255 151.685 ;
        RECT 68.855 151.640 69.145 151.685 ;
        RECT 71.975 151.640 72.265 151.685 ;
        RECT 66.965 151.500 72.265 151.640 ;
        RECT 66.965 151.455 67.255 151.500 ;
        RECT 68.855 151.455 69.145 151.500 ;
        RECT 71.975 151.455 72.265 151.500 ;
        RECT 73.440 151.640 73.760 151.700 ;
        RECT 77.085 151.640 77.375 151.685 ;
        RECT 78.975 151.640 79.265 151.685 ;
        RECT 82.095 151.640 82.385 151.685 ;
        RECT 73.440 151.500 76.890 151.640 ;
        RECT 73.440 151.440 73.760 151.500 ;
        RECT 60.560 151.300 60.880 151.360 ;
        RECT 61.955 151.300 62.245 151.345 ;
        RECT 60.560 151.160 62.245 151.300 ;
        RECT 60.560 151.100 60.880 151.160 ;
        RECT 61.955 151.115 62.245 151.160 ;
        RECT 74.820 151.100 75.140 151.360 ;
        RECT 76.750 151.300 76.890 151.500 ;
        RECT 77.085 151.500 82.385 151.640 ;
        RECT 77.085 151.455 77.375 151.500 ;
        RECT 78.975 151.455 79.265 151.500 ;
        RECT 82.095 151.455 82.385 151.500 ;
        RECT 83.650 151.300 83.790 152.180 ;
        RECT 86.320 152.120 86.640 152.180 ;
        RECT 87.240 152.120 87.560 152.380 ;
        RECT 87.720 152.320 88.010 152.365 ;
        RECT 89.555 152.320 89.845 152.365 ;
        RECT 93.135 152.320 93.425 152.365 ;
        RECT 87.720 152.180 93.425 152.320 ;
        RECT 87.720 152.135 88.010 152.180 ;
        RECT 89.555 152.135 89.845 152.180 ;
        RECT 93.135 152.135 93.425 152.180 ;
        RECT 94.215 152.160 94.505 152.475 ;
        RECT 96.455 152.320 96.745 152.365 ;
        RECT 96.070 152.180 96.745 152.320 ;
        RECT 88.620 151.780 88.940 152.040 ;
        RECT 96.070 152.025 96.210 152.180 ;
        RECT 96.455 152.135 96.745 152.180 ;
        RECT 95.995 151.795 96.285 152.025 ;
        RECT 88.125 151.640 88.415 151.685 ;
        RECT 90.015 151.640 90.305 151.685 ;
        RECT 93.135 151.640 93.425 151.685 ;
        RECT 88.125 151.500 93.425 151.640 ;
        RECT 88.125 151.455 88.415 151.500 ;
        RECT 90.015 151.455 90.305 151.500 ;
        RECT 93.135 151.455 93.425 151.500 ;
        RECT 76.750 151.160 83.790 151.300 ;
        RECT 84.940 151.100 85.260 151.360 ;
        RECT 94.140 151.300 94.460 151.360 ;
        RECT 96.915 151.300 97.205 151.345 ;
        RECT 94.140 151.160 97.205 151.300 ;
        RECT 94.140 151.100 94.460 151.160 ;
        RECT 96.915 151.115 97.205 151.160 ;
        RECT 35.190 150.480 109.250 150.960 ;
        RECT 56.830 150.280 57.120 150.325 ;
        RECT 56.830 150.140 62.170 150.280 ;
        RECT 56.830 150.095 57.120 150.140 ;
        RECT 56.385 149.940 56.675 149.985 ;
        RECT 58.275 149.940 58.565 149.985 ;
        RECT 61.395 149.940 61.685 149.985 ;
        RECT 56.385 149.800 61.685 149.940 ;
        RECT 56.385 149.755 56.675 149.800 ;
        RECT 58.275 149.755 58.565 149.800 ;
        RECT 61.395 149.755 61.685 149.800 ;
        RECT 55.515 149.600 55.805 149.645 ;
        RECT 56.880 149.600 57.200 149.660 ;
        RECT 55.515 149.460 57.200 149.600 ;
        RECT 62.030 149.600 62.170 150.140 ;
        RECT 64.240 150.080 64.560 150.340 ;
        RECT 67.920 150.280 68.240 150.340 ;
        RECT 71.140 150.280 71.460 150.340 ;
        RECT 71.615 150.280 71.905 150.325 ;
        RECT 67.920 150.140 70.910 150.280 ;
        RECT 67.920 150.080 68.240 150.140 ;
        RECT 64.330 149.600 64.470 150.080 ;
        RECT 65.160 149.940 65.480 150.000 ;
        RECT 68.855 149.940 69.145 149.985 ;
        RECT 65.160 149.800 69.145 149.940 ;
        RECT 70.770 149.940 70.910 150.140 ;
        RECT 71.140 150.140 71.905 150.280 ;
        RECT 71.140 150.080 71.460 150.140 ;
        RECT 71.615 150.095 71.905 150.140 ;
        RECT 84.020 150.280 84.340 150.340 ;
        RECT 84.495 150.280 84.785 150.325 ;
        RECT 84.020 150.140 84.785 150.280 ;
        RECT 84.020 150.080 84.340 150.140 ;
        RECT 84.495 150.095 84.785 150.140 ;
        RECT 91.380 150.080 91.700 150.340 ;
        RECT 73.440 149.940 73.760 150.000 ;
        RECT 70.770 149.800 73.760 149.940 ;
        RECT 65.160 149.740 65.480 149.800 ;
        RECT 68.855 149.755 69.145 149.800 ;
        RECT 64.715 149.600 65.005 149.645 ;
        RECT 70.695 149.600 70.985 149.645 ;
        RECT 62.030 149.460 64.010 149.600 ;
        RECT 64.330 149.460 65.005 149.600 ;
        RECT 55.515 149.415 55.805 149.460 ;
        RECT 56.880 149.400 57.200 149.460 ;
        RECT 55.980 149.260 56.270 149.305 ;
        RECT 57.815 149.260 58.105 149.305 ;
        RECT 61.395 149.260 61.685 149.305 ;
        RECT 55.980 149.120 61.685 149.260 ;
        RECT 55.980 149.075 56.270 149.120 ;
        RECT 57.815 149.075 58.105 149.120 ;
        RECT 61.395 149.075 61.685 149.120 ;
        RECT 59.175 148.920 59.825 148.965 ;
        RECT 60.560 148.920 60.880 148.980 ;
        RECT 62.475 148.965 62.765 149.280 ;
        RECT 63.870 149.260 64.010 149.460 ;
        RECT 64.715 149.415 65.005 149.460 ;
        RECT 66.860 149.460 70.985 149.600 ;
        RECT 66.860 149.260 67.000 149.460 ;
        RECT 70.695 149.415 70.985 149.460 ;
        RECT 71.230 149.305 71.370 149.800 ;
        RECT 73.440 149.740 73.760 149.800 ;
        RECT 85.860 149.940 86.180 150.000 ;
        RECT 86.335 149.940 86.625 149.985 ;
        RECT 85.860 149.800 86.625 149.940 ;
        RECT 85.860 149.740 86.180 149.800 ;
        RECT 86.335 149.755 86.625 149.800 ;
        RECT 74.820 149.600 75.140 149.660 ;
        RECT 77.135 149.600 77.425 149.645 ;
        RECT 74.820 149.460 77.425 149.600 ;
        RECT 74.820 149.400 75.140 149.460 ;
        RECT 77.135 149.415 77.425 149.460 ;
        RECT 87.255 149.600 87.545 149.645 ;
        RECT 94.140 149.600 94.460 149.660 ;
        RECT 87.255 149.460 94.460 149.600 ;
        RECT 87.255 149.415 87.545 149.460 ;
        RECT 94.140 149.400 94.460 149.460 ;
        RECT 63.870 149.120 67.000 149.260 ;
        RECT 67.935 149.260 68.225 149.305 ;
        RECT 68.395 149.260 68.685 149.305 ;
        RECT 69.775 149.260 70.065 149.305 ;
        RECT 67.935 149.120 68.685 149.260 ;
        RECT 67.935 149.075 68.225 149.120 ;
        RECT 68.395 149.075 68.685 149.120 ;
        RECT 68.930 149.120 70.065 149.260 ;
        RECT 62.475 148.920 63.065 148.965 ;
        RECT 59.175 148.780 63.065 148.920 ;
        RECT 59.175 148.735 59.825 148.780 ;
        RECT 60.560 148.720 60.880 148.780 ;
        RECT 62.775 148.735 63.065 148.780 ;
        RECT 63.320 148.920 63.640 148.980 ;
        RECT 68.930 148.920 69.070 149.120 ;
        RECT 69.775 149.075 70.065 149.120 ;
        RECT 71.155 149.075 71.445 149.305 ;
        RECT 73.440 149.260 73.760 149.320 ;
        RECT 78.055 149.260 78.345 149.305 ;
        RECT 73.440 149.120 78.345 149.260 ;
        RECT 73.440 149.060 73.760 149.120 ;
        RECT 78.055 149.075 78.345 149.120 ;
        RECT 84.940 149.060 85.260 149.320 ;
        RECT 85.875 149.075 86.165 149.305 ;
        RECT 86.320 149.260 86.640 149.320 ;
        RECT 90.935 149.260 91.225 149.305 ;
        RECT 86.320 149.120 91.225 149.260 ;
        RECT 78.500 148.920 78.820 148.980 ;
        RECT 63.320 148.780 69.070 148.920 ;
        RECT 69.390 148.780 78.820 148.920 ;
        RECT 63.320 148.720 63.640 148.780 ;
        RECT 60.100 148.580 60.420 148.640 ;
        RECT 67.000 148.580 67.320 148.640 ;
        RECT 69.390 148.580 69.530 148.780 ;
        RECT 78.500 148.720 78.820 148.780 ;
        RECT 81.720 148.920 82.040 148.980 ;
        RECT 85.950 148.920 86.090 149.075 ;
        RECT 86.320 149.060 86.640 149.120 ;
        RECT 90.935 149.075 91.225 149.120 ;
        RECT 81.720 148.780 86.090 148.920 ;
        RECT 81.720 148.720 82.040 148.780 ;
        RECT 60.100 148.440 69.530 148.580 ;
        RECT 70.680 148.580 71.000 148.640 ;
        RECT 74.375 148.580 74.665 148.625 ;
        RECT 70.680 148.440 74.665 148.580 ;
        RECT 60.100 148.380 60.420 148.440 ;
        RECT 67.000 148.380 67.320 148.440 ;
        RECT 70.680 148.380 71.000 148.440 ;
        RECT 74.375 148.395 74.665 148.440 ;
        RECT 74.820 148.580 75.140 148.640 ;
        RECT 78.975 148.580 79.265 148.625 ;
        RECT 74.820 148.440 79.265 148.580 ;
        RECT 74.820 148.380 75.140 148.440 ;
        RECT 78.975 148.395 79.265 148.440 ;
        RECT 87.255 148.580 87.545 148.625 ;
        RECT 89.080 148.580 89.400 148.640 ;
        RECT 87.255 148.440 89.400 148.580 ;
        RECT 87.255 148.395 87.545 148.440 ;
        RECT 89.080 148.380 89.400 148.440 ;
        RECT 35.190 147.760 110.030 148.240 ;
        RECT 58.735 147.560 59.025 147.605 ;
        RECT 63.320 147.560 63.640 147.620 ;
        RECT 58.735 147.420 63.640 147.560 ;
        RECT 58.735 147.375 59.025 147.420 ;
        RECT 63.320 147.360 63.640 147.420 ;
        RECT 67.460 147.560 67.780 147.620 ;
        RECT 68.395 147.560 68.685 147.605 ;
        RECT 72.075 147.560 72.365 147.605 ;
        RECT 67.460 147.420 68.685 147.560 ;
        RECT 67.460 147.360 67.780 147.420 ;
        RECT 68.395 147.375 68.685 147.420 ;
        RECT 71.690 147.420 72.365 147.560 ;
        RECT 58.260 147.220 58.580 147.280 ;
        RECT 58.260 147.080 71.370 147.220 ;
        RECT 58.260 147.020 58.580 147.080 ;
        RECT 51.820 146.680 52.140 146.940 ;
        RECT 56.435 146.880 56.725 146.925 ;
        RECT 56.435 146.740 59.410 146.880 ;
        RECT 56.435 146.695 56.725 146.740 ;
        RECT 47.680 146.340 48.000 146.600 ;
        RECT 57.340 146.340 57.660 146.600 ;
        RECT 58.260 146.340 58.580 146.600 ;
        RECT 59.270 146.540 59.410 146.740 ;
        RECT 60.100 146.680 60.420 146.940 ;
        RECT 60.575 146.880 60.865 146.925 ;
        RECT 66.080 146.880 66.400 146.940 ;
        RECT 67.935 146.880 68.225 146.925 ;
        RECT 60.575 146.740 64.010 146.880 ;
        RECT 60.575 146.695 60.865 146.740 ;
        RECT 61.020 146.540 61.340 146.600 ;
        RECT 59.270 146.400 61.340 146.540 ;
        RECT 61.020 146.340 61.340 146.400 ;
        RECT 61.480 146.540 61.800 146.600 ;
        RECT 62.415 146.540 62.705 146.585 ;
        RECT 61.480 146.400 62.705 146.540 ;
        RECT 63.870 146.540 64.010 146.740 ;
        RECT 66.080 146.740 68.225 146.880 ;
        RECT 66.080 146.680 66.400 146.740 ;
        RECT 67.935 146.695 68.225 146.740 ;
        RECT 68.380 146.880 68.700 146.940 ;
        RECT 69.315 146.880 69.605 146.925 ;
        RECT 68.380 146.740 69.605 146.880 ;
        RECT 68.380 146.680 68.700 146.740 ;
        RECT 69.315 146.695 69.605 146.740 ;
        RECT 70.680 146.680 71.000 146.940 ;
        RECT 63.870 146.400 67.000 146.540 ;
        RECT 61.480 146.340 61.800 146.400 ;
        RECT 62.415 146.355 62.705 146.400 ;
        RECT 64.700 146.200 65.020 146.260 ;
        RECT 57.430 146.060 65.020 146.200 ;
        RECT 51.360 145.660 51.680 145.920 ;
        RECT 56.420 145.860 56.740 145.920 ;
        RECT 57.430 145.905 57.570 146.060 ;
        RECT 64.700 146.000 65.020 146.060 ;
        RECT 65.160 146.200 65.480 146.260 ;
        RECT 66.095 146.200 66.385 146.245 ;
        RECT 65.160 146.060 66.385 146.200 ;
        RECT 66.860 146.200 67.000 146.400 ;
        RECT 67.460 146.340 67.780 146.600 ;
        RECT 70.220 146.540 70.540 146.600 ;
        RECT 71.230 146.540 71.370 147.080 ;
        RECT 71.690 146.925 71.830 147.420 ;
        RECT 72.075 147.375 72.365 147.420 ;
        RECT 76.675 147.560 76.965 147.605 ;
        RECT 77.580 147.560 77.900 147.620 ;
        RECT 83.100 147.560 83.420 147.620 ;
        RECT 76.675 147.420 77.900 147.560 ;
        RECT 76.675 147.375 76.965 147.420 ;
        RECT 77.580 147.360 77.900 147.420 ;
        RECT 78.130 147.420 83.420 147.560 ;
        RECT 72.995 147.220 73.285 147.265 ;
        RECT 78.130 147.220 78.270 147.420 ;
        RECT 83.100 147.360 83.420 147.420 ;
        RECT 88.620 147.560 88.940 147.620 ;
        RECT 90.015 147.560 90.305 147.605 ;
        RECT 88.620 147.420 90.305 147.560 ;
        RECT 88.620 147.360 88.940 147.420 ;
        RECT 90.015 147.375 90.305 147.420 ;
        RECT 84.495 147.220 84.785 147.265 ;
        RECT 72.995 147.080 78.270 147.220 ;
        RECT 79.970 147.080 84.785 147.220 ;
        RECT 72.995 147.035 73.285 147.080 ;
        RECT 71.615 146.695 71.905 146.925 ;
        RECT 74.835 146.880 75.125 146.925 ;
        RECT 72.610 146.740 75.125 146.880 ;
        RECT 72.610 146.540 72.750 146.740 ;
        RECT 74.835 146.695 75.125 146.740 ;
        RECT 75.280 146.680 75.600 146.940 ;
        RECT 76.215 146.695 76.505 146.925 ;
        RECT 77.595 146.880 77.885 146.925 ;
        RECT 78.040 146.880 78.360 146.940 ;
        RECT 79.970 146.925 80.110 147.080 ;
        RECT 84.495 147.035 84.785 147.080 ;
        RECT 85.415 147.220 85.705 147.265 ;
        RECT 88.175 147.220 88.465 147.265 ;
        RECT 85.415 147.080 88.465 147.220 ;
        RECT 85.415 147.035 85.705 147.080 ;
        RECT 88.175 147.035 88.465 147.080 ;
        RECT 77.595 146.740 78.360 146.880 ;
        RECT 77.595 146.695 77.885 146.740 ;
        RECT 70.220 146.400 72.750 146.540 ;
        RECT 74.360 146.540 74.680 146.600 ;
        RECT 76.290 146.540 76.430 146.695 ;
        RECT 78.040 146.680 78.360 146.740 ;
        RECT 78.515 146.880 78.805 146.925 ;
        RECT 78.515 146.740 79.650 146.880 ;
        RECT 78.515 146.695 78.805 146.740 ;
        RECT 74.360 146.400 76.430 146.540 ;
        RECT 70.220 146.340 70.540 146.400 ;
        RECT 74.360 146.340 74.680 146.400 ;
        RECT 78.960 146.340 79.280 146.600 ;
        RECT 79.510 146.540 79.650 146.740 ;
        RECT 79.895 146.695 80.185 146.925 ;
        RECT 80.815 146.880 81.105 146.925 ;
        RECT 82.180 146.880 82.500 146.940 ;
        RECT 80.815 146.740 82.500 146.880 ;
        RECT 80.815 146.695 81.105 146.740 ;
        RECT 80.890 146.540 81.030 146.695 ;
        RECT 82.180 146.680 82.500 146.740 ;
        RECT 82.640 146.680 82.960 146.940 ;
        RECT 83.100 146.680 83.420 146.940 ;
        RECT 84.955 146.880 85.245 146.925 ;
        RECT 83.650 146.740 85.245 146.880 ;
        RECT 79.510 146.400 81.030 146.540 ;
        RECT 81.275 146.540 81.565 146.585 ;
        RECT 82.730 146.540 82.870 146.680 ;
        RECT 83.650 146.540 83.790 146.740 ;
        RECT 84.955 146.695 85.245 146.740 ;
        RECT 85.860 146.680 86.180 146.940 ;
        RECT 86.320 146.880 86.640 146.940 ;
        RECT 87.255 146.880 87.545 146.925 ;
        RECT 86.320 146.740 87.545 146.880 ;
        RECT 86.320 146.680 86.640 146.740 ;
        RECT 87.255 146.695 87.545 146.740 ;
        RECT 88.635 146.695 88.925 146.925 ;
        RECT 81.275 146.400 83.790 146.540 ;
        RECT 84.020 146.540 84.340 146.600 ;
        RECT 84.495 146.540 84.785 146.585 ;
        RECT 84.020 146.400 84.785 146.540 ;
        RECT 81.275 146.355 81.565 146.400 ;
        RECT 84.020 146.340 84.340 146.400 ;
        RECT 84.495 146.355 84.785 146.400 ;
        RECT 66.860 146.060 67.690 146.200 ;
        RECT 65.160 146.000 65.480 146.060 ;
        RECT 66.095 146.015 66.385 146.060 ;
        RECT 56.895 145.860 57.185 145.905 ;
        RECT 56.420 145.720 57.185 145.860 ;
        RECT 56.420 145.660 56.740 145.720 ;
        RECT 56.895 145.675 57.185 145.720 ;
        RECT 57.355 145.675 57.645 145.905 ;
        RECT 58.260 145.860 58.580 145.920 ;
        RECT 59.655 145.860 59.945 145.905 ;
        RECT 58.260 145.720 59.945 145.860 ;
        RECT 58.260 145.660 58.580 145.720 ;
        RECT 59.655 145.675 59.945 145.720 ;
        RECT 65.620 145.660 65.940 145.920 ;
        RECT 67.000 145.660 67.320 145.920 ;
        RECT 67.550 145.860 67.690 146.060 ;
        RECT 69.760 146.000 70.080 146.260 ;
        RECT 75.755 146.200 76.045 146.245 ;
        RECT 78.055 146.200 78.345 146.245 ;
        RECT 81.720 146.200 82.040 146.260 ;
        RECT 70.310 146.060 82.040 146.200 ;
        RECT 70.310 145.860 70.450 146.060 ;
        RECT 75.755 146.015 76.045 146.060 ;
        RECT 78.055 146.015 78.345 146.060 ;
        RECT 81.720 146.000 82.040 146.060 ;
        RECT 82.655 146.200 82.945 146.245 ;
        RECT 88.710 146.200 88.850 146.695 ;
        RECT 89.080 146.680 89.400 146.940 ;
        RECT 82.655 146.060 88.850 146.200 ;
        RECT 82.655 146.015 82.945 146.060 ;
        RECT 67.550 145.720 70.450 145.860 ;
        RECT 70.680 145.860 71.000 145.920 ;
        RECT 72.995 145.860 73.285 145.905 ;
        RECT 73.440 145.860 73.760 145.920 ;
        RECT 70.680 145.720 73.760 145.860 ;
        RECT 70.680 145.660 71.000 145.720 ;
        RECT 72.995 145.675 73.285 145.720 ;
        RECT 73.440 145.660 73.760 145.720 ;
        RECT 78.500 145.860 78.820 145.920 ;
        RECT 80.815 145.860 81.105 145.905 ;
        RECT 78.500 145.720 81.105 145.860 ;
        RECT 78.500 145.660 78.820 145.720 ;
        RECT 80.815 145.675 81.105 145.720 ;
        RECT 82.180 145.860 82.500 145.920 ;
        RECT 83.560 145.860 83.880 145.920 ;
        RECT 85.860 145.860 86.180 145.920 ;
        RECT 82.180 145.720 86.180 145.860 ;
        RECT 82.180 145.660 82.500 145.720 ;
        RECT 83.560 145.660 83.880 145.720 ;
        RECT 85.860 145.660 86.180 145.720 ;
        RECT 35.190 145.040 109.250 145.520 ;
        RECT 56.435 144.840 56.725 144.885 ;
        RECT 56.880 144.840 57.200 144.900 ;
        RECT 56.435 144.700 57.200 144.840 ;
        RECT 56.435 144.655 56.725 144.700 ;
        RECT 56.880 144.640 57.200 144.700 ;
        RECT 57.340 144.840 57.660 144.900 ;
        RECT 62.860 144.840 63.180 144.900 ;
        RECT 57.340 144.700 63.180 144.840 ;
        RECT 57.340 144.640 57.660 144.700 ;
        RECT 62.860 144.640 63.180 144.700 ;
        RECT 67.460 144.840 67.780 144.900 ;
        RECT 76.200 144.840 76.520 144.900 ;
        RECT 67.460 144.700 76.520 144.840 ;
        RECT 67.460 144.640 67.780 144.700 ;
        RECT 76.200 144.640 76.520 144.700 ;
        RECT 82.655 144.840 82.945 144.885 ;
        RECT 84.480 144.840 84.800 144.900 ;
        RECT 86.320 144.840 86.640 144.900 ;
        RECT 82.655 144.700 86.640 144.840 ;
        RECT 82.655 144.655 82.945 144.700 ;
        RECT 84.480 144.640 84.800 144.700 ;
        RECT 86.320 144.640 86.640 144.700 ;
        RECT 96.455 144.840 96.745 144.885 ;
        RECT 97.820 144.840 98.140 144.900 ;
        RECT 96.455 144.700 98.140 144.840 ;
        RECT 96.455 144.655 96.745 144.700 ;
        RECT 97.820 144.640 98.140 144.700 ;
        RECT 69.760 144.500 70.080 144.560 ;
        RECT 74.820 144.500 75.140 144.560 ;
        RECT 66.860 144.360 75.140 144.500 ;
        RECT 56.420 144.160 56.740 144.220 ;
        RECT 60.560 144.160 60.880 144.220 ;
        RECT 66.860 144.160 67.000 144.360 ;
        RECT 69.760 144.300 70.080 144.360 ;
        RECT 74.820 144.300 75.140 144.360 ;
        RECT 56.420 144.020 67.000 144.160 ;
        RECT 74.910 144.020 82.410 144.160 ;
        RECT 56.420 143.960 56.740 144.020 ;
        RECT 60.560 143.960 60.880 144.020 ;
        RECT 63.795 143.820 64.085 143.865 ;
        RECT 74.360 143.820 74.680 143.880 ;
        RECT 74.910 143.865 75.050 144.020 ;
        RECT 74.835 143.820 75.125 143.865 ;
        RECT 63.795 143.680 67.000 143.820 ;
        RECT 63.795 143.635 64.085 143.680 ;
        RECT 64.700 143.280 65.020 143.540 ;
        RECT 66.860 143.480 67.000 143.680 ;
        RECT 74.360 143.680 75.125 143.820 ;
        RECT 74.360 143.620 74.680 143.680 ;
        RECT 74.835 143.635 75.125 143.680 ;
        RECT 75.280 143.820 75.600 143.880 ;
        RECT 77.120 143.820 77.440 143.880 ;
        RECT 80.800 143.820 81.120 143.880 ;
        RECT 81.720 143.820 82.040 143.880 ;
        RECT 82.270 143.865 82.410 144.020 ;
        RECT 75.280 143.680 82.040 143.820 ;
        RECT 75.280 143.620 75.600 143.680 ;
        RECT 77.120 143.620 77.440 143.680 ;
        RECT 80.800 143.620 81.120 143.680 ;
        RECT 81.720 143.620 82.040 143.680 ;
        RECT 82.195 143.635 82.485 143.865 ;
        RECT 95.980 143.620 96.300 143.880 ;
        RECT 73.440 143.480 73.760 143.540 ;
        RECT 66.860 143.340 73.760 143.480 ;
        RECT 73.440 143.280 73.760 143.340 ;
        RECT 75.755 143.480 76.045 143.525 ;
        RECT 83.100 143.480 83.420 143.540 ;
        RECT 75.755 143.340 83.420 143.480 ;
        RECT 75.755 143.295 76.045 143.340 ;
        RECT 62.860 143.140 63.180 143.200 ;
        RECT 75.830 143.140 75.970 143.295 ;
        RECT 83.100 143.280 83.420 143.340 ;
        RECT 62.860 143.000 75.970 143.140 ;
        RECT 62.860 142.940 63.180 143.000 ;
        RECT 35.190 142.320 110.030 142.800 ;
        RECT 56.880 142.120 57.200 142.180 ;
        RECT 43.170 141.980 52.050 142.120 ;
        RECT 43.170 141.780 43.310 141.980 ;
        RECT 42.710 141.640 43.310 141.780 ;
        RECT 46.295 141.780 46.945 141.825 ;
        RECT 49.895 141.780 50.185 141.825 ;
        RECT 51.360 141.780 51.680 141.840 ;
        RECT 46.295 141.640 51.680 141.780 ;
        RECT 42.710 141.485 42.850 141.640 ;
        RECT 46.295 141.595 46.945 141.640 ;
        RECT 49.595 141.595 50.185 141.640 ;
        RECT 42.635 141.255 42.925 141.485 ;
        RECT 43.100 141.440 43.390 141.485 ;
        RECT 44.935 141.440 45.225 141.485 ;
        RECT 48.515 141.440 48.805 141.485 ;
        RECT 43.100 141.300 48.805 141.440 ;
        RECT 43.100 141.255 43.390 141.300 ;
        RECT 44.935 141.255 45.225 141.300 ;
        RECT 48.515 141.255 48.805 141.300 ;
        RECT 49.595 141.280 49.885 141.595 ;
        RECT 51.360 141.580 51.680 141.640 ;
        RECT 51.910 141.780 52.050 141.980 ;
        RECT 54.670 141.980 57.200 142.120 ;
        RECT 54.670 141.840 54.810 141.980 ;
        RECT 56.880 141.920 57.200 141.980 ;
        RECT 60.575 142.120 60.865 142.165 ;
        RECT 61.480 142.120 61.800 142.180 ;
        RECT 66.080 142.120 66.400 142.180 ;
        RECT 60.575 141.980 61.800 142.120 ;
        RECT 60.575 141.935 60.865 141.980 ;
        RECT 61.480 141.920 61.800 141.980 ;
        RECT 62.490 141.980 66.400 142.120 ;
        RECT 54.580 141.780 54.900 141.840 ;
        RECT 55.960 141.825 56.280 141.840 ;
        RECT 51.910 141.640 54.900 141.780 ;
        RECT 51.910 141.485 52.050 141.640 ;
        RECT 54.580 141.580 54.900 141.640 ;
        RECT 55.495 141.780 56.280 141.825 ;
        RECT 59.095 141.780 59.385 141.825 ;
        RECT 55.495 141.640 59.385 141.780 ;
        RECT 55.495 141.595 56.280 141.640 ;
        RECT 55.960 141.580 56.280 141.595 ;
        RECT 58.795 141.595 59.385 141.640 ;
        RECT 51.835 141.255 52.125 141.485 ;
        RECT 52.300 141.440 52.590 141.485 ;
        RECT 54.135 141.440 54.425 141.485 ;
        RECT 57.715 141.440 58.005 141.485 ;
        RECT 52.300 141.300 58.005 141.440 ;
        RECT 52.300 141.255 52.590 141.300 ;
        RECT 54.135 141.255 54.425 141.300 ;
        RECT 57.715 141.255 58.005 141.300 ;
        RECT 58.795 141.280 59.085 141.595 ;
        RECT 61.020 141.580 61.340 141.840 ;
        RECT 61.110 141.440 61.250 141.580 ;
        RECT 61.480 141.440 61.800 141.500 ;
        RECT 62.490 141.485 62.630 141.980 ;
        RECT 66.080 141.920 66.400 141.980 ;
        RECT 70.680 142.120 71.000 142.180 ;
        RECT 73.455 142.120 73.745 142.165 ;
        RECT 74.820 142.120 75.140 142.180 ;
        RECT 70.680 141.980 73.745 142.120 ;
        RECT 70.680 141.920 71.000 141.980 ;
        RECT 73.455 141.935 73.745 141.980 ;
        RECT 73.990 141.980 75.140 142.120 ;
        RECT 64.715 141.780 65.005 141.825 ;
        RECT 65.160 141.780 65.480 141.840 ;
        RECT 64.715 141.640 65.480 141.780 ;
        RECT 64.715 141.595 65.005 141.640 ;
        RECT 65.160 141.580 65.480 141.640 ;
        RECT 62.415 141.440 62.705 141.485 ;
        RECT 61.110 141.300 62.705 141.440 ;
        RECT 61.480 141.240 61.800 141.300 ;
        RECT 62.415 141.255 62.705 141.300 ;
        RECT 62.860 141.240 63.180 141.500 ;
        RECT 64.255 141.440 64.545 141.485 ;
        RECT 65.620 141.440 65.940 141.500 ;
        RECT 64.255 141.300 65.940 141.440 ;
        RECT 64.255 141.255 64.545 141.300 ;
        RECT 65.620 141.240 65.940 141.300 ;
        RECT 66.095 141.255 66.385 141.485 ;
        RECT 44.015 141.100 44.305 141.145 ;
        RECT 47.680 141.100 48.000 141.160 ;
        RECT 44.015 140.960 48.000 141.100 ;
        RECT 44.015 140.915 44.305 140.960 ;
        RECT 47.680 140.900 48.000 140.960 ;
        RECT 53.215 141.100 53.505 141.145 ;
        RECT 62.950 141.100 63.090 141.240 ;
        RECT 65.160 141.100 65.480 141.160 ;
        RECT 53.215 140.960 61.710 141.100 ;
        RECT 62.950 140.960 65.480 141.100 ;
        RECT 53.215 140.915 53.505 140.960 ;
        RECT 61.570 140.805 61.710 140.960 ;
        RECT 65.160 140.900 65.480 140.960 ;
        RECT 43.505 140.760 43.795 140.805 ;
        RECT 45.395 140.760 45.685 140.805 ;
        RECT 48.515 140.760 48.805 140.805 ;
        RECT 43.505 140.620 48.805 140.760 ;
        RECT 43.505 140.575 43.795 140.620 ;
        RECT 45.395 140.575 45.685 140.620 ;
        RECT 48.515 140.575 48.805 140.620 ;
        RECT 52.705 140.760 52.995 140.805 ;
        RECT 54.595 140.760 54.885 140.805 ;
        RECT 57.715 140.760 58.005 140.805 ;
        RECT 52.705 140.620 58.005 140.760 ;
        RECT 52.705 140.575 52.995 140.620 ;
        RECT 54.595 140.575 54.885 140.620 ;
        RECT 57.715 140.575 58.005 140.620 ;
        RECT 61.495 140.575 61.785 140.805 ;
        RECT 64.240 140.760 64.560 140.820 ;
        RECT 66.170 140.760 66.310 141.255 ;
        RECT 67.000 141.240 67.320 141.500 ;
        RECT 71.155 141.440 71.445 141.485 ;
        RECT 73.440 141.440 73.760 141.500 ;
        RECT 73.990 141.485 74.130 141.980 ;
        RECT 74.820 141.920 75.140 141.980 ;
        RECT 76.200 142.120 76.520 142.180 ;
        RECT 76.200 141.980 80.110 142.120 ;
        RECT 76.200 141.920 76.520 141.980 ;
        RECT 74.375 141.780 74.665 141.825 ;
        RECT 75.280 141.780 75.600 141.840 ;
        RECT 78.960 141.780 79.280 141.840 ;
        RECT 74.375 141.640 79.280 141.780 ;
        RECT 74.375 141.595 74.665 141.640 ;
        RECT 75.280 141.580 75.600 141.640 ;
        RECT 78.960 141.580 79.280 141.640 ;
        RECT 67.550 141.300 73.760 141.440 ;
        RECT 64.240 140.620 66.310 140.760 ;
        RECT 64.240 140.560 64.560 140.620 ;
        RECT 51.375 140.420 51.665 140.465 ;
        RECT 67.550 140.420 67.690 141.300 ;
        RECT 71.155 141.255 71.445 141.300 ;
        RECT 73.440 141.240 73.760 141.300 ;
        RECT 73.915 141.255 74.205 141.485 ;
        RECT 74.835 141.255 75.125 141.485 ;
        RECT 75.755 141.440 76.045 141.485 ;
        RECT 77.120 141.440 77.440 141.500 ;
        RECT 79.970 141.485 80.110 141.980 ;
        RECT 81.275 141.935 81.565 142.165 ;
        RECT 81.350 141.780 81.490 141.935 ;
        RECT 95.980 141.920 96.300 142.180 ;
        RECT 83.345 141.780 83.635 141.825 ;
        RECT 81.350 141.640 83.635 141.780 ;
        RECT 83.345 141.595 83.635 141.640 ;
        RECT 84.480 141.580 84.800 141.840 ;
        RECT 85.875 141.780 86.165 141.825 ;
        RECT 88.635 141.780 88.925 141.825 ;
        RECT 85.875 141.640 88.925 141.780 ;
        RECT 85.875 141.595 86.165 141.640 ;
        RECT 88.635 141.595 88.925 141.640 ;
        RECT 90.915 141.780 91.565 141.825 ;
        RECT 94.515 141.780 94.805 141.825 ;
        RECT 90.915 141.640 94.805 141.780 ;
        RECT 90.915 141.595 91.565 141.640 ;
        RECT 94.215 141.595 94.805 141.640 ;
        RECT 75.755 141.300 77.440 141.440 ;
        RECT 75.755 141.255 76.045 141.300 ;
        RECT 70.220 141.100 70.540 141.160 ;
        RECT 74.910 141.100 75.050 141.255 ;
        RECT 70.220 140.960 75.050 141.100 ;
        RECT 70.220 140.900 70.540 140.960 ;
        RECT 75.830 140.760 75.970 141.255 ;
        RECT 77.120 141.240 77.440 141.300 ;
        RECT 78.515 141.440 78.805 141.485 ;
        RECT 78.515 141.300 79.650 141.440 ;
        RECT 78.515 141.255 78.805 141.300 ;
        RECT 73.070 140.620 75.970 140.760 ;
        RECT 79.510 140.760 79.650 141.300 ;
        RECT 79.895 141.255 80.185 141.485 ;
        RECT 80.800 141.440 81.120 141.500 ;
        RECT 84.020 141.440 84.340 141.500 ;
        RECT 80.800 141.300 84.340 141.440 ;
        RECT 80.800 141.240 81.120 141.300 ;
        RECT 84.020 141.240 84.340 141.300 ;
        RECT 84.940 141.240 85.260 141.500 ;
        RECT 87.720 141.440 88.010 141.485 ;
        RECT 89.555 141.440 89.845 141.485 ;
        RECT 93.135 141.440 93.425 141.485 ;
        RECT 87.720 141.300 93.425 141.440 ;
        RECT 87.720 141.255 88.010 141.300 ;
        RECT 89.555 141.255 89.845 141.300 ;
        RECT 93.135 141.255 93.425 141.300 ;
        RECT 94.215 141.440 94.505 141.595 ;
        RECT 95.520 141.440 95.840 141.500 ;
        RECT 94.215 141.300 95.840 141.440 ;
        RECT 94.215 141.280 94.505 141.300 ;
        RECT 95.520 141.240 95.840 141.300 ;
        RECT 82.640 140.900 82.960 141.160 ;
        RECT 87.240 140.900 87.560 141.160 ;
        RECT 84.940 140.760 85.260 140.820 ;
        RECT 79.510 140.620 85.260 140.760 ;
        RECT 51.375 140.280 67.690 140.420 ;
        RECT 72.535 140.420 72.825 140.465 ;
        RECT 73.070 140.420 73.210 140.620 ;
        RECT 84.940 140.560 85.260 140.620 ;
        RECT 88.125 140.760 88.415 140.805 ;
        RECT 90.015 140.760 90.305 140.805 ;
        RECT 93.135 140.760 93.425 140.805 ;
        RECT 88.125 140.620 93.425 140.760 ;
        RECT 88.125 140.575 88.415 140.620 ;
        RECT 90.015 140.575 90.305 140.620 ;
        RECT 93.135 140.575 93.425 140.620 ;
        RECT 72.535 140.280 73.210 140.420 ;
        RECT 73.440 140.420 73.760 140.480 ;
        RECT 74.360 140.420 74.680 140.480 ;
        RECT 73.440 140.280 74.680 140.420 ;
        RECT 51.375 140.235 51.665 140.280 ;
        RECT 72.535 140.235 72.825 140.280 ;
        RECT 73.440 140.220 73.760 140.280 ;
        RECT 74.360 140.220 74.680 140.280 ;
        RECT 78.960 140.220 79.280 140.480 ;
        RECT 35.190 139.600 109.250 140.080 ;
        RECT 55.960 139.200 56.280 139.460 ;
        RECT 70.220 139.400 70.540 139.460 ;
        RECT 70.695 139.400 70.985 139.445 ;
        RECT 70.220 139.260 70.985 139.400 ;
        RECT 70.220 139.200 70.540 139.260 ;
        RECT 70.695 139.215 70.985 139.260 ;
        RECT 73.900 139.400 74.220 139.460 ;
        RECT 82.640 139.400 82.960 139.460 ;
        RECT 94.155 139.400 94.445 139.445 ;
        RECT 73.900 139.260 78.270 139.400 ;
        RECT 73.900 139.200 74.220 139.260 ;
        RECT 60.575 139.060 60.865 139.105 ;
        RECT 61.480 139.060 61.800 139.120 ;
        RECT 60.575 138.920 61.800 139.060 ;
        RECT 60.575 138.875 60.865 138.920 ;
        RECT 61.480 138.860 61.800 138.920 ;
        RECT 64.240 139.060 64.560 139.120 ;
        RECT 64.240 138.920 70.910 139.060 ;
        RECT 64.240 138.860 64.560 138.920 ;
        RECT 63.335 138.720 63.625 138.765 ;
        RECT 66.095 138.720 66.385 138.765 ;
        RECT 63.335 138.580 66.385 138.720 ;
        RECT 63.335 138.535 63.625 138.580 ;
        RECT 66.095 138.535 66.385 138.580 ;
        RECT 70.770 138.720 70.910 138.920 ;
        RECT 78.130 138.720 78.270 139.260 ;
        RECT 82.640 139.260 94.445 139.400 ;
        RECT 82.640 139.200 82.960 139.260 ;
        RECT 94.155 139.215 94.445 139.260 ;
        RECT 95.520 139.200 95.840 139.460 ;
        RECT 105.195 139.400 105.485 139.445 ;
        RECT 107.480 139.400 107.800 139.460 ;
        RECT 105.195 139.260 107.800 139.400 ;
        RECT 105.195 139.215 105.485 139.260 ;
        RECT 107.480 139.200 107.800 139.260 ;
        RECT 79.435 139.060 79.725 139.105 ;
        RECT 83.560 139.060 83.880 139.120 ;
        RECT 93.695 139.060 93.985 139.105 ;
        RECT 79.435 138.920 93.985 139.060 ;
        RECT 79.435 138.875 79.725 138.920 ;
        RECT 83.560 138.860 83.880 138.920 ;
        RECT 93.695 138.875 93.985 138.920 ;
        RECT 94.615 138.720 94.905 138.765 ;
        RECT 97.820 138.720 98.140 138.780 ;
        RECT 70.770 138.580 77.350 138.720 ;
        RECT 78.130 138.580 80.570 138.720 ;
        RECT 70.770 138.440 70.910 138.580 ;
        RECT 55.500 138.180 55.820 138.440 ;
        RECT 60.100 138.180 60.420 138.440 ;
        RECT 60.560 138.380 60.880 138.440 ;
        RECT 61.035 138.380 61.325 138.425 ;
        RECT 60.560 138.240 61.325 138.380 ;
        RECT 60.560 138.180 60.880 138.240 ;
        RECT 61.035 138.195 61.325 138.240 ;
        RECT 61.495 138.380 61.785 138.425 ;
        RECT 62.415 138.380 62.705 138.425 ;
        RECT 61.495 138.240 62.705 138.380 ;
        RECT 61.495 138.195 61.785 138.240 ;
        RECT 62.415 138.195 62.705 138.240 ;
        RECT 63.795 138.380 64.085 138.425 ;
        RECT 64.240 138.380 64.560 138.440 ;
        RECT 63.795 138.240 64.560 138.380 ;
        RECT 63.795 138.195 64.085 138.240 ;
        RECT 61.110 138.040 61.250 138.195 ;
        RECT 64.240 138.180 64.560 138.240 ;
        RECT 65.160 138.180 65.480 138.440 ;
        RECT 65.620 138.180 65.940 138.440 ;
        RECT 66.540 138.380 66.860 138.440 ;
        RECT 70.680 138.425 71.000 138.440 ;
        RECT 75.830 138.425 75.970 138.580 ;
        RECT 68.855 138.380 69.145 138.425 ;
        RECT 66.540 138.240 69.145 138.380 ;
        RECT 66.540 138.180 66.860 138.240 ;
        RECT 68.855 138.195 69.145 138.240 ;
        RECT 70.680 138.195 71.135 138.425 ;
        RECT 71.615 138.195 71.905 138.425 ;
        RECT 75.755 138.195 76.045 138.425 ;
        RECT 76.675 138.195 76.965 138.425 ;
        RECT 77.210 138.390 77.350 138.580 ;
        RECT 80.430 138.425 80.570 138.580 ;
        RECT 94.615 138.580 98.140 138.720 ;
        RECT 94.615 138.535 94.905 138.580 ;
        RECT 97.820 138.520 98.140 138.580 ;
        RECT 77.595 138.390 77.885 138.425 ;
        RECT 77.210 138.250 77.885 138.390 ;
        RECT 77.595 138.195 77.885 138.250 ;
        RECT 78.975 138.195 79.265 138.425 ;
        RECT 80.355 138.195 80.645 138.425 ;
        RECT 92.775 138.195 93.065 138.425 ;
        RECT 70.680 138.180 71.000 138.195 ;
        RECT 65.710 138.040 65.850 138.180 ;
        RECT 71.690 138.040 71.830 138.195 ;
        RECT 76.750 138.040 76.890 138.195 ;
        RECT 79.050 138.040 79.190 138.195 ;
        RECT 79.420 138.040 79.740 138.100 ;
        RECT 61.110 137.900 65.850 138.040 ;
        RECT 69.390 137.900 79.740 138.040 ;
        RECT 69.390 137.760 69.530 137.900 ;
        RECT 79.420 137.840 79.740 137.900 ;
        RECT 82.180 138.040 82.500 138.100 ;
        RECT 89.555 138.040 89.845 138.085 ;
        RECT 82.180 137.900 89.845 138.040 ;
        RECT 92.850 138.040 92.990 138.195 ;
        RECT 93.220 138.180 93.540 138.440 ;
        RECT 95.060 138.180 95.380 138.440 ;
        RECT 95.980 138.380 96.300 138.440 ;
        RECT 104.735 138.380 105.025 138.425 ;
        RECT 95.980 138.240 105.025 138.380 ;
        RECT 95.980 138.180 96.300 138.240 ;
        RECT 104.735 138.195 105.025 138.240 ;
        RECT 96.070 138.040 96.210 138.180 ;
        RECT 92.850 137.900 96.210 138.040 ;
        RECT 82.180 137.840 82.500 137.900 ;
        RECT 89.555 137.855 89.845 137.900 ;
        RECT 59.180 137.500 59.500 137.760 ;
        RECT 64.715 137.700 65.005 137.745 ;
        RECT 67.000 137.700 67.320 137.760 ;
        RECT 69.300 137.700 69.620 137.760 ;
        RECT 64.715 137.560 69.620 137.700 ;
        RECT 64.715 137.515 65.005 137.560 ;
        RECT 67.000 137.500 67.320 137.560 ;
        RECT 69.300 137.500 69.620 137.560 ;
        RECT 76.215 137.700 76.505 137.745 ;
        RECT 78.040 137.700 78.360 137.760 ;
        RECT 84.940 137.700 85.260 137.760 ;
        RECT 76.215 137.560 85.260 137.700 ;
        RECT 76.215 137.515 76.505 137.560 ;
        RECT 78.040 137.500 78.360 137.560 ;
        RECT 84.940 137.500 85.260 137.560 ;
        RECT 86.795 137.700 87.085 137.745 ;
        RECT 87.240 137.700 87.560 137.760 ;
        RECT 86.795 137.560 87.560 137.700 ;
        RECT 86.795 137.515 87.085 137.560 ;
        RECT 87.240 137.500 87.560 137.560 ;
        RECT 35.190 136.880 110.030 137.360 ;
        RECT 60.575 136.680 60.865 136.725 ;
        RECT 63.780 136.680 64.100 136.740 ;
        RECT 66.540 136.680 66.860 136.740 ;
        RECT 60.575 136.540 66.860 136.680 ;
        RECT 60.575 136.495 60.865 136.540 ;
        RECT 63.780 136.480 64.100 136.540 ;
        RECT 66.540 136.480 66.860 136.540 ;
        RECT 77.580 136.680 77.900 136.740 ;
        RECT 93.220 136.680 93.540 136.740 ;
        RECT 77.580 136.540 93.540 136.680 ;
        RECT 77.580 136.480 77.900 136.540 ;
        RECT 53.200 136.340 53.520 136.400 ;
        RECT 54.580 136.340 54.900 136.400 ;
        RECT 51.910 136.200 54.900 136.340 ;
        RECT 51.910 136.045 52.050 136.200 ;
        RECT 53.200 136.140 53.520 136.200 ;
        RECT 54.580 136.140 54.900 136.200 ;
        RECT 55.495 136.340 56.145 136.385 ;
        RECT 59.095 136.340 59.385 136.385 ;
        RECT 61.955 136.340 62.245 136.385 ;
        RECT 55.495 136.200 62.245 136.340 ;
        RECT 55.495 136.155 56.145 136.200 ;
        RECT 58.795 136.155 59.385 136.200 ;
        RECT 61.955 136.155 62.245 136.200 ;
        RECT 73.455 136.340 73.745 136.385 ;
        RECT 74.375 136.340 74.665 136.385 ;
        RECT 73.455 136.200 74.665 136.340 ;
        RECT 73.455 136.155 73.745 136.200 ;
        RECT 74.375 136.155 74.665 136.200 ;
        RECT 75.740 136.340 76.060 136.400 ;
        RECT 78.960 136.340 79.280 136.400 ;
        RECT 79.435 136.340 79.725 136.385 ;
        RECT 75.740 136.200 79.725 136.340 ;
        RECT 51.835 135.815 52.125 136.045 ;
        RECT 52.300 136.000 52.590 136.045 ;
        RECT 54.135 136.000 54.425 136.045 ;
        RECT 57.715 136.000 58.005 136.045 ;
        RECT 52.300 135.860 58.005 136.000 ;
        RECT 52.300 135.815 52.590 135.860 ;
        RECT 54.135 135.815 54.425 135.860 ;
        RECT 57.715 135.815 58.005 135.860 ;
        RECT 58.795 135.840 59.085 136.155 ;
        RECT 75.740 136.140 76.060 136.200 ;
        RECT 78.960 136.140 79.280 136.200 ;
        RECT 79.435 136.155 79.725 136.200 ;
        RECT 81.720 136.340 82.040 136.400 ;
        RECT 84.110 136.385 84.250 136.540 ;
        RECT 93.220 136.480 93.540 136.540 ;
        RECT 95.980 136.480 96.300 136.740 ;
        RECT 82.885 136.340 83.175 136.385 ;
        RECT 81.720 136.200 83.175 136.340 ;
        RECT 81.720 136.140 82.040 136.200 ;
        RECT 82.885 136.155 83.175 136.200 ;
        RECT 84.035 136.155 84.325 136.385 ;
        RECT 85.415 136.340 85.705 136.385 ;
        RECT 88.635 136.340 88.925 136.385 ;
        RECT 85.415 136.200 88.925 136.340 ;
        RECT 85.415 136.155 85.705 136.200 ;
        RECT 88.635 136.155 88.925 136.200 ;
        RECT 90.000 136.340 90.320 136.400 ;
        RECT 90.915 136.340 91.565 136.385 ;
        RECT 94.515 136.340 94.805 136.385 ;
        RECT 90.000 136.200 94.805 136.340 ;
        RECT 90.000 136.140 90.320 136.200 ;
        RECT 90.915 136.155 91.565 136.200 ;
        RECT 94.215 136.155 94.805 136.200 ;
        RECT 62.415 136.000 62.705 136.045 ;
        RECT 66.095 136.000 66.385 136.045 ;
        RECT 67.460 136.000 67.780 136.060 ;
        RECT 68.840 136.000 69.160 136.060 ;
        RECT 62.415 135.860 69.160 136.000 ;
        RECT 62.415 135.815 62.705 135.860 ;
        RECT 66.095 135.815 66.385 135.860 ;
        RECT 67.460 135.800 67.780 135.860 ;
        RECT 68.840 135.800 69.160 135.860 ;
        RECT 73.915 135.815 74.205 136.045 ;
        RECT 53.215 135.660 53.505 135.705 ;
        RECT 59.180 135.660 59.500 135.720 ;
        RECT 53.215 135.520 59.500 135.660 ;
        RECT 53.215 135.475 53.505 135.520 ;
        RECT 59.180 135.460 59.500 135.520 ;
        RECT 69.300 135.660 69.620 135.720 ;
        RECT 70.235 135.660 70.525 135.705 ;
        RECT 69.300 135.520 70.525 135.660 ;
        RECT 73.990 135.660 74.130 135.815 ;
        RECT 75.280 135.800 75.600 136.060 ;
        RECT 77.580 135.800 77.900 136.060 ;
        RECT 78.040 135.800 78.360 136.060 ;
        RECT 79.880 135.990 80.200 136.060 ;
        RECT 80.815 136.000 81.105 136.045 ;
        RECT 80.430 135.990 81.105 136.000 ;
        RECT 79.880 135.860 81.105 135.990 ;
        RECT 79.880 135.850 80.570 135.860 ;
        RECT 79.880 135.800 80.200 135.850 ;
        RECT 80.815 135.815 81.105 135.860 ;
        RECT 82.180 135.800 82.500 136.060 ;
        RECT 83.560 135.800 83.880 136.060 ;
        RECT 84.495 136.000 84.785 136.045 ;
        RECT 84.940 136.000 85.260 136.060 ;
        RECT 84.495 135.860 85.260 136.000 ;
        RECT 84.495 135.815 84.785 135.860 ;
        RECT 84.940 135.800 85.260 135.860 ;
        RECT 87.720 136.000 88.010 136.045 ;
        RECT 89.555 136.000 89.845 136.045 ;
        RECT 93.135 136.000 93.425 136.045 ;
        RECT 87.720 135.860 93.425 136.000 ;
        RECT 87.720 135.815 88.010 135.860 ;
        RECT 89.555 135.815 89.845 135.860 ;
        RECT 93.135 135.815 93.425 135.860 ;
        RECT 94.215 135.840 94.505 136.155 ;
        RECT 74.820 135.660 75.140 135.720 ;
        RECT 77.670 135.660 77.810 135.800 ;
        RECT 73.990 135.520 77.810 135.660 ;
        RECT 69.300 135.460 69.620 135.520 ;
        RECT 70.235 135.475 70.525 135.520 ;
        RECT 74.820 135.460 75.140 135.520 ;
        RECT 78.975 135.475 79.265 135.705 ;
        RECT 80.355 135.660 80.645 135.705 ;
        RECT 82.640 135.660 82.960 135.720 ;
        RECT 80.355 135.520 82.960 135.660 ;
        RECT 80.355 135.475 80.645 135.520 ;
        RECT 52.705 135.320 52.995 135.365 ;
        RECT 54.595 135.320 54.885 135.365 ;
        RECT 57.715 135.320 58.005 135.365 ;
        RECT 52.705 135.180 58.005 135.320 ;
        RECT 52.705 135.135 52.995 135.180 ;
        RECT 54.595 135.135 54.885 135.180 ;
        RECT 57.715 135.135 58.005 135.180 ;
        RECT 66.555 135.320 66.845 135.365 ;
        RECT 67.000 135.320 67.320 135.380 ;
        RECT 66.555 135.180 67.320 135.320 ;
        RECT 79.050 135.320 79.190 135.475 ;
        RECT 82.640 135.460 82.960 135.520 ;
        RECT 83.650 135.320 83.790 135.800 ;
        RECT 87.240 135.460 87.560 135.720 ;
        RECT 79.050 135.180 83.790 135.320 ;
        RECT 88.125 135.320 88.415 135.365 ;
        RECT 90.015 135.320 90.305 135.365 ;
        RECT 93.135 135.320 93.425 135.365 ;
        RECT 88.125 135.180 93.425 135.320 ;
        RECT 66.555 135.135 66.845 135.180 ;
        RECT 67.000 135.120 67.320 135.180 ;
        RECT 88.125 135.135 88.415 135.180 ;
        RECT 90.015 135.135 90.305 135.180 ;
        RECT 93.135 135.135 93.425 135.180 ;
        RECT 76.200 134.780 76.520 135.040 ;
        RECT 78.500 134.780 78.820 135.040 ;
        RECT 79.420 134.780 79.740 135.040 ;
        RECT 81.720 134.780 82.040 135.040 ;
        RECT 35.190 134.160 109.250 134.640 ;
        RECT 79.880 133.960 80.200 134.020 ;
        RECT 77.210 133.820 80.200 133.960 ;
        RECT 61.960 133.620 62.250 133.665 ;
        RECT 63.820 133.620 64.110 133.665 ;
        RECT 66.600 133.620 66.890 133.665 ;
        RECT 61.960 133.480 66.890 133.620 ;
        RECT 61.960 133.435 62.250 133.480 ;
        RECT 63.820 133.435 64.110 133.480 ;
        RECT 66.600 133.435 66.890 133.480 ;
        RECT 53.200 133.280 53.520 133.340 ;
        RECT 70.680 133.325 71.000 133.340 ;
        RECT 77.210 133.325 77.350 133.820 ;
        RECT 79.880 133.760 80.200 133.820 ;
        RECT 82.640 133.960 82.960 134.020 ;
        RECT 84.020 133.960 84.340 134.020 ;
        RECT 86.795 133.960 87.085 134.005 ;
        RECT 82.640 133.820 87.085 133.960 ;
        RECT 82.640 133.760 82.960 133.820 ;
        RECT 84.020 133.760 84.340 133.820 ;
        RECT 86.795 133.775 87.085 133.820 ;
        RECT 90.000 133.760 90.320 134.020 ;
        RECT 78.515 133.620 78.805 133.665 ;
        RECT 80.355 133.620 80.645 133.665 ;
        RECT 83.115 133.620 83.405 133.665 ;
        RECT 78.515 133.480 83.405 133.620 ;
        RECT 78.515 133.435 78.805 133.480 ;
        RECT 80.355 133.435 80.645 133.480 ;
        RECT 83.115 133.435 83.405 133.480 ;
        RECT 61.495 133.280 61.785 133.325 ;
        RECT 70.465 133.280 71.000 133.325 ;
        RECT 77.135 133.280 77.425 133.325 ;
        RECT 87.240 133.280 87.560 133.340 ;
        RECT 53.200 133.140 61.785 133.280 ;
        RECT 70.245 133.140 77.425 133.280 ;
        RECT 53.200 133.080 53.520 133.140 ;
        RECT 61.495 133.095 61.785 133.140 ;
        RECT 70.465 133.095 71.000 133.140 ;
        RECT 77.135 133.095 77.425 133.140 ;
        RECT 78.130 133.140 87.560 133.280 ;
        RECT 70.680 133.080 71.000 133.095 ;
        RECT 78.130 133.000 78.270 133.140 ;
        RECT 87.240 133.080 87.560 133.140 ;
        RECT 63.335 132.940 63.625 132.985 ;
        RECT 63.780 132.940 64.100 133.000 ;
        RECT 66.600 132.940 66.890 132.985 ;
        RECT 63.335 132.800 64.100 132.940 ;
        RECT 63.335 132.755 63.625 132.800 ;
        RECT 63.780 132.740 64.100 132.800 ;
        RECT 64.355 132.800 66.890 132.940 ;
        RECT 64.355 132.645 64.570 132.800 ;
        RECT 66.600 132.755 66.890 132.800 ;
        RECT 67.460 132.940 67.780 133.000 ;
        RECT 73.455 132.940 73.745 132.985 ;
        RECT 67.460 132.800 77.350 132.940 ;
        RECT 67.460 132.740 67.780 132.800 ;
        RECT 73.455 132.755 73.745 132.800 ;
        RECT 62.420 132.600 62.710 132.645 ;
        RECT 64.280 132.600 64.570 132.645 ;
        RECT 62.420 132.460 64.570 132.600 ;
        RECT 62.420 132.415 62.710 132.460 ;
        RECT 64.280 132.415 64.570 132.460 ;
        RECT 65.200 132.600 65.490 132.645 ;
        RECT 67.000 132.600 67.320 132.660 ;
        RECT 68.460 132.600 68.750 132.645 ;
        RECT 65.200 132.460 68.750 132.600 ;
        RECT 65.200 132.415 65.490 132.460 ;
        RECT 67.000 132.400 67.320 132.460 ;
        RECT 68.460 132.415 68.750 132.460 ;
        RECT 72.995 132.260 73.285 132.305 ;
        RECT 73.440 132.260 73.760 132.320 ;
        RECT 72.995 132.120 73.760 132.260 ;
        RECT 72.995 132.075 73.285 132.120 ;
        RECT 73.440 132.060 73.760 132.120 ;
        RECT 74.360 132.060 74.680 132.320 ;
        RECT 77.210 132.260 77.350 132.800 ;
        RECT 78.040 132.740 78.360 133.000 ;
        RECT 78.500 132.940 78.820 133.000 ;
        RECT 79.895 132.940 80.185 132.985 ;
        RECT 83.135 132.940 83.425 132.985 ;
        RECT 78.500 132.800 80.185 132.940 ;
        RECT 78.500 132.740 78.820 132.800 ;
        RECT 79.895 132.755 80.185 132.800 ;
        RECT 80.890 132.800 83.425 132.940 ;
        RECT 80.890 132.645 81.105 132.800 ;
        RECT 83.135 132.755 83.425 132.800 ;
        RECT 84.020 132.940 84.340 133.000 ;
        RECT 89.555 132.940 89.845 132.985 ;
        RECT 95.060 132.940 95.380 133.000 ;
        RECT 84.020 132.800 95.380 132.940 ;
        RECT 84.020 132.740 84.340 132.800 ;
        RECT 89.555 132.755 89.845 132.800 ;
        RECT 95.060 132.740 95.380 132.800 ;
        RECT 78.975 132.600 79.265 132.645 ;
        RECT 80.815 132.600 81.105 132.645 ;
        RECT 78.975 132.460 81.105 132.600 ;
        RECT 78.975 132.415 79.265 132.460 ;
        RECT 80.815 132.415 81.105 132.460 ;
        RECT 81.735 132.600 82.025 132.645 ;
        RECT 83.560 132.600 83.880 132.660 ;
        RECT 84.955 132.600 85.245 132.645 ;
        RECT 81.735 132.460 85.245 132.600 ;
        RECT 81.735 132.415 82.025 132.460 ;
        RECT 83.560 132.400 83.880 132.460 ;
        RECT 84.955 132.415 85.245 132.460 ;
        RECT 84.020 132.260 84.340 132.320 ;
        RECT 77.210 132.120 84.340 132.260 ;
        RECT 84.020 132.060 84.340 132.120 ;
        RECT 35.190 131.440 110.030 131.920 ;
        RECT 63.780 131.040 64.100 131.300 ;
        RECT 83.560 131.040 83.880 131.300 ;
        RECT 71.155 130.900 71.445 130.945 ;
        RECT 73.440 130.900 73.760 130.960 ;
        RECT 74.375 130.900 74.665 130.945 ;
        RECT 71.155 130.760 74.665 130.900 ;
        RECT 71.155 130.715 71.445 130.760 ;
        RECT 73.440 130.700 73.760 130.760 ;
        RECT 74.375 130.715 74.665 130.760 ;
        RECT 75.295 130.900 75.585 130.945 ;
        RECT 77.135 130.900 77.425 130.945 ;
        RECT 75.295 130.760 77.425 130.900 ;
        RECT 75.295 130.715 75.585 130.760 ;
        RECT 77.135 130.715 77.425 130.760 ;
        RECT 72.975 130.560 73.265 130.605 ;
        RECT 75.295 130.560 75.510 130.715 ;
        RECT 72.975 130.420 75.510 130.560 ;
        RECT 72.975 130.375 73.265 130.420 ;
        RECT 76.200 130.360 76.520 130.620 ;
        RECT 78.040 130.360 78.360 130.620 ;
        RECT 84.020 130.360 84.340 130.620 ;
        RECT 67.000 130.020 67.320 130.280 ;
        RECT 72.995 129.880 73.285 129.925 ;
        RECT 75.755 129.880 76.045 129.925 ;
        RECT 77.595 129.880 77.885 129.925 ;
        RECT 72.995 129.740 77.885 129.880 ;
        RECT 72.995 129.695 73.285 129.740 ;
        RECT 75.755 129.695 76.045 129.740 ;
        RECT 77.595 129.695 77.885 129.740 ;
        RECT 69.300 129.340 69.620 129.600 ;
        RECT 35.190 128.720 109.250 129.200 ;
        RECT 63.795 128.180 64.085 128.225 ;
        RECT 67.000 128.180 67.320 128.240 ;
        RECT 63.795 128.040 67.320 128.180 ;
        RECT 63.795 127.995 64.085 128.040 ;
        RECT 67.000 127.980 67.320 128.040 ;
        RECT 74.360 127.840 74.680 127.900 ;
        RECT 64.790 127.700 74.680 127.840 ;
        RECT 64.790 127.545 64.930 127.700 ;
        RECT 74.360 127.640 74.680 127.700 ;
        RECT 64.715 127.315 65.005 127.545 ;
        RECT 65.620 127.300 65.940 127.560 ;
        RECT 66.095 127.500 66.385 127.545 ;
        RECT 69.300 127.500 69.620 127.560 ;
        RECT 66.095 127.360 69.620 127.500 ;
        RECT 66.095 127.315 66.385 127.360 ;
        RECT 69.300 127.300 69.620 127.360 ;
        RECT 35.190 126.000 110.030 126.480 ;
        RECT 35.190 123.280 109.250 123.760 ;
        RECT 35.190 120.560 110.030 121.040 ;
        RECT 35.190 117.840 109.250 118.320 ;
        RECT 35.190 115.120 110.030 115.600 ;
        RECT 35.190 112.400 109.250 112.880 ;
        RECT 35.190 109.680 110.030 110.160 ;
        RECT 35.190 106.960 109.250 107.440 ;
        RECT 35.190 104.240 110.030 104.720 ;
        RECT 35.190 101.520 109.250 102.000 ;
        RECT 35.190 98.800 110.030 99.280 ;
        RECT 35.190 96.080 109.250 96.560 ;
        RECT 35.190 93.360 110.030 93.840 ;
        RECT 35.190 90.640 109.250 91.120 ;
        RECT 35.190 87.920 110.030 88.400 ;
        RECT 35.190 85.200 109.250 85.680 ;
        RECT 75.280 84.800 75.600 85.060 ;
        RECT 74.820 83.440 75.140 83.700 ;
        RECT 35.190 82.480 110.030 82.960 ;
        RECT 72.520 82.280 72.840 82.340 ;
        RECT 74.820 82.280 75.140 82.340 ;
        RECT 72.520 82.140 75.140 82.280 ;
        RECT 72.520 82.080 72.840 82.140 ;
        RECT 74.820 82.080 75.140 82.140 ;
        RECT 105.060 79.000 137.720 79.010 ;
        RECT 105.010 77.210 137.720 79.000 ;
        RECT 105.010 77.200 110.680 77.210 ;
        RECT 105.010 77.190 107.880 77.200 ;
        RECT 20.000 76.550 22.000 77.050 ;
        RECT 20.000 76.250 37.050 76.550 ;
        RECT 20.000 75.955 22.400 76.250 ;
        RECT 20.000 75.820 22.870 75.955 ;
        RECT 23.050 75.820 23.550 75.900 ;
        RECT 28.800 75.820 29.300 75.900 ;
        RECT 20.000 75.590 23.780 75.820 ;
        RECT 20.000 75.455 22.870 75.590 ;
        RECT 23.050 75.510 23.550 75.590 ;
        RECT 20.000 74.400 22.400 75.455 ;
        RECT 22.800 75.030 23.300 75.110 ;
        RECT 22.780 74.800 23.780 75.030 ;
        RECT 23.920 75.010 24.220 75.610 ;
        RECT 25.935 75.010 26.235 75.610 ;
        RECT 26.375 75.590 36.375 75.820 ;
        RECT 28.800 75.510 29.300 75.590 ;
        RECT 29.800 75.030 30.800 75.110 ;
        RECT 26.375 74.800 36.375 75.030 ;
        RECT 22.800 74.720 23.300 74.800 ;
        RECT 29.800 74.720 30.800 74.800 ;
        RECT 36.750 74.400 37.050 76.250 ;
        RECT 20.000 74.100 37.050 74.400 ;
        RECT 20.000 35.000 22.000 74.100 ;
        RECT 37.200 73.300 39.200 77.050 ;
        RECT 22.150 73.000 39.200 73.300 ;
        RECT 22.150 69.750 22.450 73.000 ;
        RECT 22.800 72.690 23.300 72.770 ;
        RECT 28.800 72.690 29.300 72.770 ;
        RECT 22.730 72.460 23.730 72.690 ;
        RECT 22.800 72.380 23.300 72.460 ;
        RECT 22.730 71.900 23.230 71.980 ;
        RECT 22.730 71.670 23.730 71.900 ;
        RECT 23.900 71.880 24.200 72.480 ;
        RECT 25.950 71.880 26.250 72.480 ;
        RECT 26.420 72.460 36.420 72.690 ;
        RECT 28.800 72.380 29.300 72.460 ;
        RECT 29.800 71.900 30.800 71.980 ;
        RECT 22.730 71.590 23.230 71.670 ;
        RECT 22.730 71.110 23.230 71.190 ;
        RECT 22.730 70.880 23.730 71.110 ;
        RECT 23.900 71.090 24.200 71.690 ;
        RECT 25.950 71.090 26.250 71.690 ;
        RECT 26.420 71.670 36.420 71.900 ;
        RECT 29.800 71.585 30.800 71.670 ;
        RECT 28.800 71.110 29.300 71.190 ;
        RECT 22.730 70.800 23.230 70.880 ;
        RECT 22.730 70.320 23.230 70.400 ;
        RECT 22.730 70.090 23.730 70.320 ;
        RECT 23.900 70.300 24.200 70.900 ;
        RECT 25.950 70.300 26.250 70.900 ;
        RECT 26.420 70.880 36.420 71.110 ;
        RECT 28.800 70.800 29.300 70.880 ;
        RECT 29.800 70.320 30.800 70.400 ;
        RECT 26.420 70.090 36.420 70.320 ;
        RECT 22.730 70.010 23.230 70.090 ;
        RECT 29.800 70.010 30.800 70.090 ;
        RECT 36.700 69.750 39.200 73.000 ;
        RECT 40.000 71.050 104.800 73.050 ;
        RECT 40.000 71.000 41.050 71.050 ;
        RECT 22.150 69.450 39.200 69.750 ;
        RECT 37.200 35.000 39.200 69.450 ;
        RECT 40.350 57.150 40.950 71.000 ;
        RECT 48.500 70.710 49.100 70.740 ;
        RECT 53.140 70.710 53.740 70.740 ;
        RECT 60.030 70.710 60.630 70.740 ;
        RECT 66.920 70.710 67.520 70.740 ;
        RECT 73.810 70.710 74.410 70.740 ;
        RECT 80.700 70.710 81.300 70.740 ;
        RECT 87.590 70.710 88.190 70.740 ;
        RECT 48.300 70.480 50.800 70.710 ;
        RECT 51.440 70.480 57.690 70.710 ;
        RECT 58.330 70.480 64.580 70.710 ;
        RECT 65.220 70.480 71.470 70.710 ;
        RECT 72.110 70.480 78.360 70.710 ;
        RECT 79.000 70.480 85.250 70.710 ;
        RECT 85.890 70.480 88.390 70.710 ;
        RECT 48.500 70.450 49.100 70.480 ;
        RECT 53.140 70.450 53.740 70.480 ;
        RECT 60.030 70.450 60.630 70.480 ;
        RECT 66.920 70.450 67.520 70.480 ;
        RECT 73.810 70.450 74.410 70.480 ;
        RECT 80.700 70.450 81.300 70.480 ;
        RECT 87.590 70.450 88.190 70.480 ;
        RECT 47.865 70.370 48.095 70.430 ;
        RECT 47.750 69.530 48.200 70.370 ;
        RECT 47.865 69.470 48.095 69.530 ;
        RECT 51.005 69.470 51.235 70.430 ;
        RECT 57.895 69.470 58.125 70.430 ;
        RECT 64.785 69.470 65.015 70.430 ;
        RECT 71.675 69.470 71.905 70.430 ;
        RECT 78.565 69.470 78.795 70.430 ;
        RECT 85.455 69.470 85.685 70.430 ;
        RECT 88.595 70.370 88.825 70.430 ;
        RECT 88.500 69.530 88.950 70.370 ;
        RECT 88.595 69.470 88.825 69.530 ;
        RECT 48.500 69.420 49.100 69.450 ;
        RECT 55.390 69.420 55.990 69.450 ;
        RECT 62.280 69.420 62.880 69.450 ;
        RECT 69.170 69.420 69.770 69.450 ;
        RECT 76.060 69.420 76.660 69.450 ;
        RECT 82.950 69.420 83.550 69.450 ;
        RECT 87.590 69.420 88.190 69.450 ;
        RECT 48.300 69.190 50.800 69.420 ;
        RECT 51.440 69.190 57.690 69.420 ;
        RECT 58.330 69.190 64.580 69.420 ;
        RECT 65.220 69.190 71.470 69.420 ;
        RECT 72.110 69.190 78.360 69.420 ;
        RECT 79.000 69.190 85.250 69.420 ;
        RECT 85.890 69.190 88.390 69.420 ;
        RECT 48.500 69.160 49.100 69.190 ;
        RECT 55.390 69.160 55.990 69.190 ;
        RECT 62.280 69.160 62.880 69.190 ;
        RECT 69.170 69.160 69.770 69.190 ;
        RECT 76.060 69.160 76.660 69.190 ;
        RECT 82.950 69.160 83.550 69.190 ;
        RECT 87.590 69.160 88.190 69.190 ;
        RECT 47.865 69.080 48.095 69.140 ;
        RECT 47.750 68.240 48.200 69.080 ;
        RECT 47.865 68.180 48.095 68.240 ;
        RECT 51.005 68.180 51.235 69.140 ;
        RECT 57.895 68.180 58.125 69.140 ;
        RECT 64.785 68.180 65.015 69.140 ;
        RECT 71.675 68.180 71.905 69.140 ;
        RECT 78.565 68.180 78.795 69.140 ;
        RECT 85.455 68.180 85.685 69.140 ;
        RECT 88.595 69.080 88.825 69.140 ;
        RECT 88.500 68.240 88.950 69.080 ;
        RECT 88.595 68.180 88.825 68.240 ;
        RECT 48.500 68.130 49.100 68.160 ;
        RECT 53.140 68.130 53.740 68.160 ;
        RECT 60.030 68.130 60.630 68.160 ;
        RECT 66.920 68.130 67.520 68.160 ;
        RECT 73.805 68.130 74.405 68.160 ;
        RECT 80.700 68.130 81.300 68.160 ;
        RECT 87.590 68.130 88.190 68.160 ;
        RECT 48.300 67.900 50.800 68.130 ;
        RECT 51.440 67.900 57.690 68.130 ;
        RECT 58.330 67.900 64.580 68.130 ;
        RECT 65.220 67.900 71.470 68.130 ;
        RECT 72.110 67.900 78.360 68.130 ;
        RECT 79.000 67.900 85.250 68.130 ;
        RECT 85.890 67.900 88.390 68.130 ;
        RECT 48.500 67.870 49.100 67.900 ;
        RECT 53.140 67.870 53.740 67.900 ;
        RECT 60.030 67.870 60.630 67.900 ;
        RECT 66.920 67.870 67.520 67.900 ;
        RECT 73.805 67.870 74.405 67.900 ;
        RECT 80.700 67.870 81.300 67.900 ;
        RECT 87.590 67.870 88.190 67.900 ;
        RECT 47.865 67.790 48.095 67.850 ;
        RECT 47.750 66.950 48.200 67.790 ;
        RECT 47.865 66.890 48.095 66.950 ;
        RECT 51.005 66.890 51.235 67.850 ;
        RECT 57.895 66.890 58.125 67.850 ;
        RECT 64.785 66.890 65.015 67.850 ;
        RECT 71.675 66.890 71.905 67.850 ;
        RECT 78.565 66.890 78.795 67.850 ;
        RECT 85.455 66.890 85.685 67.850 ;
        RECT 88.595 67.790 88.825 67.850 ;
        RECT 88.500 66.950 88.950 67.790 ;
        RECT 88.595 66.890 88.825 66.950 ;
        RECT 48.500 66.840 49.100 66.870 ;
        RECT 55.390 66.840 55.990 66.870 ;
        RECT 62.280 66.840 62.880 66.870 ;
        RECT 69.170 66.840 69.770 66.870 ;
        RECT 76.060 66.840 76.660 66.870 ;
        RECT 82.950 66.840 83.550 66.870 ;
        RECT 87.590 66.840 88.190 66.870 ;
        RECT 48.300 66.610 50.800 66.840 ;
        RECT 51.440 66.610 57.690 66.840 ;
        RECT 58.330 66.610 64.580 66.840 ;
        RECT 65.220 66.610 71.470 66.840 ;
        RECT 72.110 66.610 78.360 66.840 ;
        RECT 79.000 66.610 85.250 66.840 ;
        RECT 85.890 66.610 88.390 66.840 ;
        RECT 48.500 66.580 49.100 66.610 ;
        RECT 55.390 66.580 55.990 66.610 ;
        RECT 62.280 66.580 62.880 66.610 ;
        RECT 69.170 66.580 69.770 66.610 ;
        RECT 76.060 66.580 76.660 66.610 ;
        RECT 82.950 66.580 83.550 66.610 ;
        RECT 87.590 66.580 88.190 66.610 ;
        RECT 47.865 66.500 48.095 66.560 ;
        RECT 47.750 65.660 48.200 66.500 ;
        RECT 47.865 65.600 48.095 65.660 ;
        RECT 51.005 65.600 51.235 66.560 ;
        RECT 57.895 65.600 58.125 66.560 ;
        RECT 64.785 65.600 65.015 66.560 ;
        RECT 71.675 65.600 71.905 66.560 ;
        RECT 78.565 65.600 78.795 66.560 ;
        RECT 85.455 65.600 85.685 66.560 ;
        RECT 88.595 66.500 88.825 66.560 ;
        RECT 88.500 65.660 88.950 66.500 ;
        RECT 95.750 66.350 96.350 71.050 ;
        RECT 100.100 70.640 100.700 70.670 ;
        RECT 97.800 69.810 98.200 70.450 ;
        RECT 98.340 70.410 101.340 70.640 ;
        RECT 100.100 70.380 100.700 70.410 ;
        RECT 98.700 69.850 99.300 69.880 ;
        RECT 98.340 69.620 101.340 69.850 ;
        RECT 98.700 69.590 99.300 69.620 ;
        RECT 100.100 69.180 100.700 69.210 ;
        RECT 98.750 68.200 99.150 69.050 ;
        RECT 99.300 68.950 102.300 69.180 ;
        RECT 100.100 68.920 100.700 68.950 ;
        RECT 100.400 68.390 101.000 68.420 ;
        RECT 99.300 68.160 102.300 68.390 ;
        RECT 100.400 68.130 101.000 68.160 ;
        RECT 103.850 66.350 104.450 71.050 ;
        RECT 95.750 65.750 104.450 66.350 ;
        RECT 88.595 65.600 88.825 65.660 ;
        RECT 48.500 65.550 49.100 65.580 ;
        RECT 53.140 65.550 53.740 65.580 ;
        RECT 60.030 65.550 60.630 65.580 ;
        RECT 66.920 65.550 67.520 65.580 ;
        RECT 73.810 65.550 74.410 65.580 ;
        RECT 80.700 65.550 81.300 65.580 ;
        RECT 87.590 65.550 88.190 65.580 ;
        RECT 48.300 65.320 50.800 65.550 ;
        RECT 51.440 65.320 57.690 65.550 ;
        RECT 58.330 65.320 64.580 65.550 ;
        RECT 65.220 65.320 71.470 65.550 ;
        RECT 72.110 65.320 78.360 65.550 ;
        RECT 79.000 65.320 85.250 65.550 ;
        RECT 85.890 65.320 88.390 65.550 ;
        RECT 48.500 65.290 49.100 65.320 ;
        RECT 53.140 65.290 53.740 65.320 ;
        RECT 60.030 65.290 60.630 65.320 ;
        RECT 66.920 65.290 67.520 65.320 ;
        RECT 73.810 65.290 74.410 65.320 ;
        RECT 80.700 65.290 81.300 65.320 ;
        RECT 87.590 65.290 88.190 65.320 ;
        RECT 47.865 65.210 48.095 65.270 ;
        RECT 47.750 64.370 48.200 65.210 ;
        RECT 47.865 64.310 48.095 64.370 ;
        RECT 51.005 64.310 51.235 65.270 ;
        RECT 57.895 64.310 58.125 65.270 ;
        RECT 64.785 64.310 65.015 65.270 ;
        RECT 71.675 64.310 71.905 65.270 ;
        RECT 78.565 64.310 78.795 65.270 ;
        RECT 85.455 64.310 85.685 65.270 ;
        RECT 88.595 65.210 88.825 65.270 ;
        RECT 88.500 64.370 88.950 65.210 ;
        RECT 88.595 64.310 88.825 64.370 ;
        RECT 48.500 64.260 49.100 64.290 ;
        RECT 55.390 64.260 55.990 64.290 ;
        RECT 62.280 64.260 62.880 64.290 ;
        RECT 69.170 64.260 69.770 64.290 ;
        RECT 76.060 64.260 76.660 64.290 ;
        RECT 82.950 64.260 83.550 64.290 ;
        RECT 87.590 64.260 88.190 64.290 ;
        RECT 48.300 64.030 50.800 64.260 ;
        RECT 51.440 64.030 57.690 64.260 ;
        RECT 58.330 64.030 64.580 64.260 ;
        RECT 65.220 64.030 71.470 64.260 ;
        RECT 72.110 64.030 78.360 64.260 ;
        RECT 79.000 64.030 85.250 64.260 ;
        RECT 85.890 64.030 88.390 64.260 ;
        RECT 48.500 64.000 49.100 64.030 ;
        RECT 55.390 64.000 55.990 64.030 ;
        RECT 62.280 64.000 62.880 64.030 ;
        RECT 69.170 64.000 69.770 64.030 ;
        RECT 76.060 64.000 76.660 64.030 ;
        RECT 82.950 64.000 83.550 64.030 ;
        RECT 87.590 64.000 88.190 64.030 ;
        RECT 47.865 63.920 48.095 63.980 ;
        RECT 47.750 63.080 48.200 63.920 ;
        RECT 47.865 63.020 48.095 63.080 ;
        RECT 51.005 63.020 51.235 63.980 ;
        RECT 57.895 63.020 58.125 63.980 ;
        RECT 64.785 63.020 65.015 63.980 ;
        RECT 71.675 63.020 71.905 63.980 ;
        RECT 78.565 63.020 78.795 63.980 ;
        RECT 85.455 63.020 85.685 63.980 ;
        RECT 88.595 63.920 88.825 63.980 ;
        RECT 88.500 63.080 88.950 63.920 ;
        RECT 88.595 63.020 88.825 63.080 ;
        RECT 48.500 62.970 49.100 63.000 ;
        RECT 53.140 62.970 53.740 63.000 ;
        RECT 60.030 62.970 60.630 63.000 ;
        RECT 66.920 62.970 67.520 63.000 ;
        RECT 73.810 62.970 74.410 63.000 ;
        RECT 80.700 62.970 81.300 63.000 ;
        RECT 87.590 62.970 88.190 63.000 ;
        RECT 48.300 62.740 50.800 62.970 ;
        RECT 51.440 62.740 57.690 62.970 ;
        RECT 58.330 62.740 64.580 62.970 ;
        RECT 65.220 62.740 71.470 62.970 ;
        RECT 72.110 62.740 78.360 62.970 ;
        RECT 79.000 62.740 85.250 62.970 ;
        RECT 85.890 62.740 88.390 62.970 ;
        RECT 48.500 62.710 49.100 62.740 ;
        RECT 53.140 62.710 53.740 62.740 ;
        RECT 60.030 62.710 60.630 62.740 ;
        RECT 66.920 62.710 67.520 62.740 ;
        RECT 73.810 62.710 74.410 62.740 ;
        RECT 80.700 62.710 81.300 62.740 ;
        RECT 87.590 62.710 88.190 62.740 ;
        RECT 47.865 62.630 48.095 62.690 ;
        RECT 47.750 61.790 48.200 62.630 ;
        RECT 47.865 61.730 48.095 61.790 ;
        RECT 51.005 61.730 51.235 62.690 ;
        RECT 57.895 61.730 58.125 62.690 ;
        RECT 64.785 61.730 65.015 62.690 ;
        RECT 71.675 61.730 71.905 62.690 ;
        RECT 78.565 61.730 78.795 62.690 ;
        RECT 85.455 61.730 85.685 62.690 ;
        RECT 88.595 62.630 88.825 62.690 ;
        RECT 88.500 61.790 88.950 62.630 ;
        RECT 88.595 61.730 88.825 61.790 ;
        RECT 48.500 61.680 49.100 61.710 ;
        RECT 55.390 61.680 55.990 61.710 ;
        RECT 62.280 61.680 62.880 61.710 ;
        RECT 69.170 61.680 69.770 61.710 ;
        RECT 76.060 61.680 76.660 61.710 ;
        RECT 82.950 61.680 83.550 61.710 ;
        RECT 87.590 61.680 88.190 61.710 ;
        RECT 48.300 61.450 50.800 61.680 ;
        RECT 51.440 61.450 57.690 61.680 ;
        RECT 58.330 61.450 64.580 61.680 ;
        RECT 65.220 61.450 71.470 61.680 ;
        RECT 72.110 61.450 78.360 61.680 ;
        RECT 79.000 61.450 85.250 61.680 ;
        RECT 85.890 61.450 88.390 61.680 ;
        RECT 48.500 61.420 49.100 61.450 ;
        RECT 55.390 61.420 55.990 61.450 ;
        RECT 62.280 61.420 62.880 61.450 ;
        RECT 69.170 61.420 69.770 61.450 ;
        RECT 76.060 61.420 76.660 61.450 ;
        RECT 82.950 61.420 83.550 61.450 ;
        RECT 87.590 61.420 88.190 61.450 ;
        RECT 47.865 61.340 48.095 61.400 ;
        RECT 47.750 60.500 48.200 61.340 ;
        RECT 47.865 60.440 48.095 60.500 ;
        RECT 51.005 60.440 51.235 61.400 ;
        RECT 57.895 60.440 58.125 61.400 ;
        RECT 64.785 60.440 65.015 61.400 ;
        RECT 71.675 60.440 71.905 61.400 ;
        RECT 78.565 60.440 78.795 61.400 ;
        RECT 85.455 60.440 85.685 61.400 ;
        RECT 88.595 61.340 88.825 61.400 ;
        RECT 88.500 60.500 88.950 61.340 ;
        RECT 88.595 60.440 88.825 60.500 ;
        RECT 48.500 60.390 49.100 60.420 ;
        RECT 53.140 60.390 53.740 60.420 ;
        RECT 60.025 60.390 60.625 60.420 ;
        RECT 66.920 60.390 67.520 60.420 ;
        RECT 73.810 60.390 74.410 60.415 ;
        RECT 80.700 60.390 81.300 60.420 ;
        RECT 87.590 60.390 88.190 60.420 ;
        RECT 48.300 60.160 50.800 60.390 ;
        RECT 51.440 60.160 57.690 60.390 ;
        RECT 58.330 60.160 64.580 60.390 ;
        RECT 65.220 60.160 71.470 60.390 ;
        RECT 72.110 60.160 78.360 60.390 ;
        RECT 79.000 60.160 85.250 60.390 ;
        RECT 85.890 60.160 88.390 60.390 ;
        RECT 48.500 60.130 49.100 60.160 ;
        RECT 53.140 60.130 53.740 60.160 ;
        RECT 60.025 60.130 60.625 60.160 ;
        RECT 66.920 60.130 67.520 60.160 ;
        RECT 73.810 60.125 74.410 60.160 ;
        RECT 80.700 60.130 81.300 60.160 ;
        RECT 87.590 60.130 88.190 60.160 ;
        RECT 95.750 57.150 96.350 65.750 ;
        RECT 40.350 56.550 96.350 57.150 ;
        RECT 40.350 42.800 40.950 56.550 ;
        RECT 47.550 56.230 48.150 56.260 ;
        RECT 88.550 56.230 89.150 56.260 ;
        RECT 41.600 56.000 67.035 56.230 ;
        RECT 47.550 55.970 48.150 56.000 ;
        RECT 41.165 54.990 41.395 55.950 ;
        RECT 66.805 54.990 67.035 56.000 ;
        RECT 69.665 56.000 95.100 56.230 ;
        RECT 69.665 54.990 69.895 56.000 ;
        RECT 88.550 55.970 89.150 56.000 ;
        RECT 95.305 54.990 95.535 55.950 ;
        RECT 47.550 54.940 48.150 54.970 ;
        RECT 88.550 54.940 89.150 54.970 ;
        RECT 41.600 54.710 66.600 54.940 ;
        RECT 70.100 54.710 95.100 54.940 ;
        RECT 47.550 54.680 48.150 54.710 ;
        RECT 88.550 54.680 89.150 54.710 ;
        RECT 41.165 53.700 41.395 54.660 ;
        RECT 66.805 54.430 67.035 54.660 ;
        RECT 66.805 53.930 68.150 54.430 ;
        RECT 53.800 53.650 54.400 53.680 ;
        RECT 41.600 53.420 66.600 53.650 ;
        RECT 53.800 53.390 54.400 53.420 ;
        RECT 41.165 52.410 41.395 53.370 ;
        RECT 66.805 52.410 67.035 53.930 ;
        RECT 69.665 53.140 69.895 54.660 ;
        RECT 95.305 53.700 95.535 54.660 ;
        RECT 82.300 53.650 82.900 53.680 ;
        RECT 70.100 53.420 95.100 53.650 ;
        RECT 82.300 53.390 82.900 53.420 ;
        RECT 68.550 52.640 69.895 53.140 ;
        RECT 69.665 52.410 69.895 52.640 ;
        RECT 95.305 52.410 95.535 53.370 ;
        RECT 47.550 52.360 48.150 52.390 ;
        RECT 88.550 52.360 89.150 52.390 ;
        RECT 41.600 52.130 66.600 52.360 ;
        RECT 70.100 52.130 95.100 52.360 ;
        RECT 47.550 52.100 48.150 52.130 ;
        RECT 88.550 52.100 89.150 52.130 ;
        RECT 41.165 51.120 41.395 52.080 ;
        RECT 66.805 51.850 67.035 52.080 ;
        RECT 66.805 51.350 69.150 51.850 ;
        RECT 60.050 51.070 60.650 51.100 ;
        RECT 41.600 50.840 66.600 51.070 ;
        RECT 60.050 50.810 60.650 50.840 ;
        RECT 41.165 49.830 41.395 50.790 ;
        RECT 66.805 49.830 67.035 51.350 ;
        RECT 69.665 50.560 69.895 52.080 ;
        RECT 95.305 51.120 95.535 52.080 ;
        RECT 76.050 51.070 76.650 51.100 ;
        RECT 70.100 50.840 95.100 51.070 ;
        RECT 76.050 50.810 76.650 50.840 ;
        RECT 67.550 50.060 69.895 50.560 ;
        RECT 69.665 49.830 69.895 50.060 ;
        RECT 95.305 49.830 95.535 50.790 ;
        RECT 47.550 49.780 48.150 49.810 ;
        RECT 88.550 49.780 89.150 49.810 ;
        RECT 41.600 49.550 66.600 49.780 ;
        RECT 70.100 49.550 95.100 49.780 ;
        RECT 47.550 49.520 48.150 49.550 ;
        RECT 88.550 49.520 89.150 49.550 ;
        RECT 41.165 48.540 41.395 49.500 ;
        RECT 66.805 49.270 67.035 49.500 ;
        RECT 66.805 48.770 69.150 49.270 ;
        RECT 60.050 48.490 60.650 48.520 ;
        RECT 41.600 48.260 66.600 48.490 ;
        RECT 60.050 48.230 60.650 48.260 ;
        RECT 41.165 47.250 41.395 48.210 ;
        RECT 66.805 47.250 67.035 48.770 ;
        RECT 69.665 47.980 69.895 49.500 ;
        RECT 95.305 48.540 95.535 49.500 ;
        RECT 76.050 48.490 76.650 48.520 ;
        RECT 70.100 48.260 95.100 48.490 ;
        RECT 76.050 48.230 76.650 48.260 ;
        RECT 67.550 47.480 69.895 47.980 ;
        RECT 69.665 47.250 69.895 47.480 ;
        RECT 95.305 47.250 95.535 48.210 ;
        RECT 47.550 47.200 48.150 47.230 ;
        RECT 88.550 47.200 89.150 47.230 ;
        RECT 41.600 46.970 66.600 47.200 ;
        RECT 70.100 46.970 95.100 47.200 ;
        RECT 47.550 46.940 48.150 46.970 ;
        RECT 88.550 46.940 89.150 46.970 ;
        RECT 41.165 45.960 41.395 46.920 ;
        RECT 66.805 46.690 67.035 46.920 ;
        RECT 66.805 46.190 68.150 46.690 ;
        RECT 53.800 45.910 54.400 45.940 ;
        RECT 41.600 45.680 66.600 45.910 ;
        RECT 53.800 45.650 54.400 45.680 ;
        RECT 41.165 44.670 41.395 45.630 ;
        RECT 66.805 44.670 67.035 46.190 ;
        RECT 69.665 45.400 69.895 46.920 ;
        RECT 95.305 45.960 95.535 46.920 ;
        RECT 82.300 45.910 82.900 45.940 ;
        RECT 70.100 45.680 95.100 45.910 ;
        RECT 82.300 45.650 82.900 45.680 ;
        RECT 68.550 44.900 69.895 45.400 ;
        RECT 69.665 44.670 69.895 44.900 ;
        RECT 95.305 44.670 95.535 45.630 ;
        RECT 47.550 44.620 48.150 44.650 ;
        RECT 88.550 44.620 89.150 44.650 ;
        RECT 41.600 44.390 66.600 44.620 ;
        RECT 70.100 44.390 95.100 44.620 ;
        RECT 47.550 44.360 48.150 44.390 ;
        RECT 88.550 44.360 89.150 44.390 ;
        RECT 41.165 43.380 41.395 44.340 ;
        RECT 47.550 43.330 48.150 43.360 ;
        RECT 66.805 43.330 67.035 44.340 ;
        RECT 41.600 43.100 67.035 43.330 ;
        RECT 69.665 43.330 69.895 44.340 ;
        RECT 95.305 43.380 95.535 44.340 ;
        RECT 88.550 43.330 89.150 43.360 ;
        RECT 69.665 43.100 95.100 43.330 ;
        RECT 47.550 43.070 48.150 43.100 ;
        RECT 88.550 43.070 89.150 43.100 ;
        RECT 95.750 42.800 96.350 56.550 ;
        RECT 40.350 42.200 96.350 42.800 ;
        RECT 97.150 64.350 104.800 64.950 ;
        RECT 97.150 62.450 97.700 64.350 ;
        RECT 98.650 63.700 99.350 63.730 ;
        RECT 100.350 63.700 101.050 63.730 ;
        RECT 97.850 62.850 98.250 63.600 ;
        RECT 98.390 63.470 100.130 63.700 ;
        RECT 100.290 63.470 101.290 63.700 ;
        RECT 98.650 63.440 99.350 63.470 ;
        RECT 99.900 62.960 100.130 63.470 ;
        RECT 100.350 63.440 101.050 63.470 ;
        RECT 98.390 62.800 99.390 62.910 ;
        RECT 100.290 62.800 101.290 62.910 ;
        RECT 98.390 62.680 104.100 62.800 ;
        RECT 97.150 41.400 97.750 62.450 ;
        RECT 98.400 62.300 104.100 62.680 ;
        RECT 104.250 61.850 104.800 64.350 ;
        RECT 98.560 60.550 99.520 60.780 ;
        RECT 99.850 60.550 100.810 60.780 ;
        RECT 101.140 60.550 102.100 60.780 ;
        RECT 102.430 60.550 103.390 60.780 ;
        RECT 98.280 49.250 98.510 60.390 ;
        RECT 99.570 59.950 99.800 60.390 ;
        RECT 99.490 59.450 99.880 59.950 ;
        RECT 98.200 48.750 98.590 49.250 ;
        RECT 98.280 42.890 98.510 48.750 ;
        RECT 99.570 42.890 99.800 59.450 ;
        RECT 100.860 49.250 101.090 60.390 ;
        RECT 102.150 59.950 102.380 60.390 ;
        RECT 102.070 59.450 102.460 59.950 ;
        RECT 100.780 48.750 101.170 49.250 ;
        RECT 100.860 42.890 101.090 48.750 ;
        RECT 102.150 42.890 102.380 59.450 ;
        RECT 103.440 49.250 103.670 60.390 ;
        RECT 103.360 48.750 103.750 49.250 ;
        RECT 103.440 42.890 103.670 48.750 ;
        RECT 98.550 42.400 99.550 42.750 ;
        RECT 99.850 42.400 100.850 42.750 ;
        RECT 101.150 42.730 102.150 42.750 ;
        RECT 102.450 42.730 103.450 42.750 ;
        RECT 101.140 42.500 102.150 42.730 ;
        RECT 102.430 42.500 103.450 42.730 ;
        RECT 101.150 42.400 102.150 42.500 ;
        RECT 102.450 42.400 103.450 42.500 ;
        RECT 40.350 40.800 97.750 41.400 ;
        RECT 40.350 37.000 40.950 40.800 ;
        RECT 45.675 40.290 46.280 40.320 ;
        RECT 52.225 40.290 52.830 40.320 ;
        RECT 61.775 40.290 62.380 40.320 ;
        RECT 71.325 40.290 71.930 40.320 ;
        RECT 80.875 40.290 81.480 40.325 ;
        RECT 90.425 40.290 91.030 40.320 ;
        RECT 44.475 40.060 48.975 40.290 ;
        RECT 49.525 40.060 58.525 40.290 ;
        RECT 59.075 40.060 68.075 40.290 ;
        RECT 68.625 40.060 77.625 40.290 ;
        RECT 78.175 40.060 87.175 40.290 ;
        RECT 87.725 40.060 92.225 40.290 ;
        RECT 45.675 40.030 46.280 40.060 ;
        RECT 52.225 40.030 52.830 40.060 ;
        RECT 61.775 40.030 62.380 40.060 ;
        RECT 71.325 40.030 71.930 40.060 ;
        RECT 80.875 40.035 81.480 40.060 ;
        RECT 90.425 40.030 91.030 40.060 ;
        RECT 44.085 39.900 44.315 40.010 ;
        RECT 44.000 39.150 44.400 39.900 ;
        RECT 44.085 39.050 44.315 39.150 ;
        RECT 49.135 39.050 49.365 40.010 ;
        RECT 58.685 39.050 58.915 40.010 ;
        RECT 68.235 39.050 68.465 40.010 ;
        RECT 77.785 39.050 78.015 40.010 ;
        RECT 87.335 39.050 87.565 40.010 ;
        RECT 92.385 39.900 92.615 40.010 ;
        RECT 92.300 39.150 92.700 39.900 ;
        RECT 92.385 39.050 92.615 39.150 ;
        RECT 45.675 39.000 46.280 39.030 ;
        RECT 55.225 39.000 55.825 39.030 ;
        RECT 64.775 39.000 65.375 39.030 ;
        RECT 74.320 39.000 74.930 39.030 ;
        RECT 83.870 39.000 84.480 39.030 ;
        RECT 90.425 39.000 91.030 39.030 ;
        RECT 44.475 38.770 48.975 39.000 ;
        RECT 49.525 38.770 58.525 39.000 ;
        RECT 59.075 38.770 68.075 39.000 ;
        RECT 68.625 38.770 77.625 39.000 ;
        RECT 78.175 38.770 87.175 39.000 ;
        RECT 87.725 38.770 92.225 39.000 ;
        RECT 45.675 38.740 46.280 38.770 ;
        RECT 55.225 38.740 55.825 38.770 ;
        RECT 64.775 38.740 65.375 38.770 ;
        RECT 74.320 38.740 74.930 38.770 ;
        RECT 83.870 38.740 84.480 38.770 ;
        RECT 90.425 38.740 91.030 38.770 ;
        RECT 44.085 38.600 44.315 38.720 ;
        RECT 44.000 37.850 44.400 38.600 ;
        RECT 44.085 37.760 44.315 37.850 ;
        RECT 49.135 37.760 49.365 38.720 ;
        RECT 58.685 37.760 58.915 38.720 ;
        RECT 68.235 37.760 68.465 38.720 ;
        RECT 77.785 37.760 78.015 38.720 ;
        RECT 87.335 37.760 87.565 38.720 ;
        RECT 92.385 38.600 92.615 38.720 ;
        RECT 92.300 37.850 92.700 38.600 ;
        RECT 92.385 37.760 92.615 37.850 ;
        RECT 45.675 37.710 46.280 37.740 ;
        RECT 52.225 37.710 52.830 37.740 ;
        RECT 61.775 37.710 62.380 37.740 ;
        RECT 71.325 37.710 71.930 37.740 ;
        RECT 80.875 37.710 81.480 37.740 ;
        RECT 90.425 37.710 91.030 37.740 ;
        RECT 44.475 37.480 48.975 37.710 ;
        RECT 49.525 37.480 58.525 37.710 ;
        RECT 59.075 37.480 68.075 37.710 ;
        RECT 68.625 37.480 77.625 37.710 ;
        RECT 78.175 37.480 87.175 37.710 ;
        RECT 87.725 37.480 92.225 37.710 ;
        RECT 45.675 37.450 46.280 37.480 ;
        RECT 52.225 37.450 52.830 37.480 ;
        RECT 61.775 37.450 62.380 37.480 ;
        RECT 71.325 37.450 71.930 37.480 ;
        RECT 80.875 37.450 81.480 37.480 ;
        RECT 90.425 37.450 91.030 37.480 ;
        RECT 104.200 37.000 104.800 61.850 ;
        RECT 107.380 60.790 107.610 77.190 ;
        RECT 108.090 60.790 108.480 76.800 ;
        RECT 108.960 60.790 109.190 77.200 ;
        RECT 109.670 60.790 110.060 76.790 ;
        RECT 111.080 60.800 111.310 77.210 ;
        RECT 111.790 60.800 112.180 76.810 ;
        RECT 112.660 60.800 112.890 77.210 ;
        RECT 113.370 60.800 113.760 76.800 ;
        RECT 114.790 60.800 115.020 77.210 ;
        RECT 115.500 60.800 115.890 76.810 ;
        RECT 116.370 60.800 116.600 77.210 ;
        RECT 117.080 60.800 117.470 76.800 ;
        RECT 118.500 60.800 118.730 77.210 ;
        RECT 119.210 60.800 119.600 76.810 ;
        RECT 120.080 60.800 120.310 77.210 ;
        RECT 120.790 60.800 121.180 76.800 ;
        RECT 122.210 60.800 122.440 77.210 ;
        RECT 122.920 60.800 123.310 76.810 ;
        RECT 123.790 60.800 124.020 77.210 ;
        RECT 124.500 60.800 124.890 76.800 ;
        RECT 125.920 60.800 126.150 77.210 ;
        RECT 126.630 60.800 127.020 76.810 ;
        RECT 127.500 60.800 127.730 77.210 ;
        RECT 128.210 60.800 128.600 76.800 ;
        RECT 129.630 60.800 129.860 77.210 ;
        RECT 130.340 60.800 130.730 76.810 ;
        RECT 131.210 60.800 131.440 77.210 ;
        RECT 131.920 60.800 132.310 76.800 ;
        RECT 133.340 60.800 133.570 77.210 ;
        RECT 134.050 60.800 134.440 76.810 ;
        RECT 134.920 60.800 135.150 77.210 ;
        RECT 135.630 60.800 136.020 76.800 ;
        RECT 107.660 59.590 108.120 60.590 ;
        RECT 108.450 59.590 108.910 60.590 ;
        RECT 109.240 59.590 109.700 60.590 ;
        RECT 107.660 59.310 109.700 59.590 ;
        RECT 111.360 59.600 111.820 60.600 ;
        RECT 112.150 59.600 112.610 60.600 ;
        RECT 112.940 59.600 113.400 60.600 ;
        RECT 107.660 58.875 109.705 59.310 ;
        RECT 107.660 58.590 109.700 58.875 ;
        RECT 107.660 57.590 108.120 58.590 ;
        RECT 108.450 57.590 108.910 58.590 ;
        RECT 109.240 57.590 109.700 58.590 ;
        RECT 111.360 58.600 113.400 59.600 ;
        RECT 111.360 57.600 111.820 58.600 ;
        RECT 112.150 57.600 112.610 58.600 ;
        RECT 112.940 57.600 113.400 58.600 ;
        RECT 115.070 59.600 115.530 60.600 ;
        RECT 115.860 59.600 116.320 60.600 ;
        RECT 116.650 59.600 117.110 60.600 ;
        RECT 115.070 58.600 117.110 59.600 ;
        RECT 115.070 57.600 115.530 58.600 ;
        RECT 115.860 57.600 116.320 58.600 ;
        RECT 116.650 57.600 117.110 58.600 ;
        RECT 118.780 59.600 119.240 60.600 ;
        RECT 119.570 59.600 120.030 60.600 ;
        RECT 120.360 59.600 120.820 60.600 ;
        RECT 118.780 58.600 120.820 59.600 ;
        RECT 118.780 57.600 119.240 58.600 ;
        RECT 119.570 57.600 120.030 58.600 ;
        RECT 120.360 57.600 120.820 58.600 ;
        RECT 122.490 59.600 122.950 60.600 ;
        RECT 123.280 59.600 123.740 60.600 ;
        RECT 124.070 59.600 124.530 60.600 ;
        RECT 122.490 58.600 124.530 59.600 ;
        RECT 122.490 57.600 122.950 58.600 ;
        RECT 123.280 57.600 123.740 58.600 ;
        RECT 124.070 57.600 124.530 58.600 ;
        RECT 126.200 59.600 126.660 60.600 ;
        RECT 126.990 59.600 127.450 60.600 ;
        RECT 127.780 59.600 128.240 60.600 ;
        RECT 126.200 58.600 128.240 59.600 ;
        RECT 126.200 57.600 126.660 58.600 ;
        RECT 126.990 57.600 127.450 58.600 ;
        RECT 127.780 57.600 128.240 58.600 ;
        RECT 129.910 59.600 130.370 60.600 ;
        RECT 130.700 59.600 131.160 60.600 ;
        RECT 131.490 59.600 131.950 60.600 ;
        RECT 129.910 58.600 131.950 59.600 ;
        RECT 129.910 57.600 130.370 58.600 ;
        RECT 130.700 57.600 131.160 58.600 ;
        RECT 131.490 57.600 131.950 58.600 ;
        RECT 133.620 59.600 134.080 60.600 ;
        RECT 134.410 59.600 134.870 60.600 ;
        RECT 135.200 59.600 135.660 60.600 ;
        RECT 133.620 58.600 135.660 59.600 ;
        RECT 133.620 57.600 134.080 58.600 ;
        RECT 134.410 57.600 134.870 58.600 ;
        RECT 135.200 57.600 135.660 58.600 ;
        RECT 107.380 50.030 107.610 57.430 ;
        RECT 108.090 50.430 108.480 57.430 ;
        RECT 108.960 50.030 109.190 57.430 ;
        RECT 109.670 50.430 110.060 57.430 ;
        RECT 111.080 50.030 111.310 57.440 ;
        RECT 111.790 50.440 112.180 57.440 ;
        RECT 112.660 50.030 112.890 57.440 ;
        RECT 113.370 50.440 113.760 57.440 ;
        RECT 114.790 50.030 115.020 57.440 ;
        RECT 115.500 50.440 115.890 57.440 ;
        RECT 116.370 50.030 116.600 57.440 ;
        RECT 117.080 50.440 117.470 57.440 ;
        RECT 118.500 50.030 118.730 57.440 ;
        RECT 119.210 50.440 119.600 57.440 ;
        RECT 120.080 50.030 120.310 57.440 ;
        RECT 120.790 50.440 121.180 57.440 ;
        RECT 122.210 50.030 122.440 57.440 ;
        RECT 122.920 50.440 123.310 57.440 ;
        RECT 123.790 50.030 124.020 57.440 ;
        RECT 124.500 50.440 124.890 57.440 ;
        RECT 125.920 50.030 126.150 57.440 ;
        RECT 126.630 50.440 127.020 57.440 ;
        RECT 127.500 50.030 127.730 57.440 ;
        RECT 128.210 50.440 128.600 57.440 ;
        RECT 129.630 50.030 129.860 57.440 ;
        RECT 130.340 50.440 130.730 57.440 ;
        RECT 131.210 50.030 131.440 57.440 ;
        RECT 131.920 50.440 132.310 57.440 ;
        RECT 133.340 50.030 133.570 57.440 ;
        RECT 134.050 50.440 134.440 57.440 ;
        RECT 134.920 50.030 135.150 57.440 ;
        RECT 135.630 50.440 136.020 57.440 ;
        RECT 105.080 50.020 136.640 50.030 ;
        RECT 105.030 48.820 137.720 50.020 ;
        RECT 105.080 48.020 106.210 48.820 ;
        RECT 105.080 46.810 107.670 48.020 ;
        RECT 110.340 46.990 111.440 47.990 ;
        RECT 113.840 47.000 114.940 48.000 ;
        RECT 117.330 47.010 118.440 48.000 ;
        RECT 117.380 47.000 118.380 47.010 ;
        RECT 120.870 47.000 121.970 48.000 ;
        RECT 124.360 47.010 125.480 48.020 ;
        RECT 127.860 47.010 128.960 48.020 ;
        RECT 132.810 48.010 134.570 48.020 ;
        RECT 40.000 35.000 104.800 37.000 ;
        RECT 105.090 44.850 107.670 46.810 ;
        RECT 108.240 44.850 110.000 46.960 ;
        RECT 110.580 44.850 111.170 46.990 ;
        RECT 111.760 46.960 113.500 46.980 ;
        RECT 111.750 44.870 113.510 46.960 ;
        RECT 111.750 44.855 113.520 44.870 ;
        RECT 105.090 35.580 106.490 44.850 ;
        RECT 109.400 39.120 110.000 44.850 ;
        RECT 111.760 44.840 113.520 44.855 ;
        RECT 114.070 44.840 114.690 47.000 ;
        RECT 115.260 44.855 117.060 46.960 ;
        RECT 117.580 44.870 118.190 47.000 ;
        RECT 117.600 44.855 118.190 44.870 ;
        RECT 118.760 44.860 120.530 46.980 ;
        RECT 118.770 44.855 119.360 44.860 ;
        RECT 115.270 44.840 117.060 44.855 ;
        RECT 109.400 38.520 112.340 39.120 ;
        RECT 107.070 35.860 108.830 37.970 ;
        RECT 109.410 37.960 110.000 37.965 ;
        RECT 110.580 37.960 111.170 37.965 ;
        RECT 109.410 35.860 111.180 37.960 ;
        RECT 111.730 35.860 112.340 38.520 ;
        RECT 112.930 39.090 113.520 44.840 ;
        RECT 116.420 39.160 117.060 44.840 ;
        RECT 112.930 39.065 115.865 39.090 ;
        RECT 112.930 38.500 115.870 39.065 ;
        RECT 116.420 38.520 119.390 39.160 ;
        RECT 119.930 39.120 120.530 44.860 ;
        RECT 121.110 44.850 121.710 47.000 ;
        RECT 122.280 44.855 124.040 46.960 ;
        RECT 122.290 44.850 124.040 44.855 ;
        RECT 124.620 44.850 125.210 47.010 ;
        RECT 125.780 46.960 127.540 46.970 ;
        RECT 125.780 44.850 127.550 46.960 ;
        RECT 128.130 44.850 128.720 47.010 ;
        RECT 131.360 47.000 132.470 48.010 ;
        RECT 129.280 44.850 131.060 46.970 ;
        RECT 131.640 44.850 132.230 47.000 ;
        RECT 132.760 44.850 134.610 48.010 ;
        RECT 134.890 47.010 135.990 48.010 ;
        RECT 135.150 44.850 135.740 47.010 ;
        RECT 123.430 39.120 124.040 44.850 ;
        RECT 126.930 39.120 127.550 44.850 ;
        RECT 130.430 39.150 131.060 44.850 ;
        RECT 119.930 38.520 122.870 39.120 ;
        RECT 109.420 35.850 111.180 35.860 ;
        RECT 112.900 35.830 114.680 37.980 ;
        RECT 115.260 35.860 115.870 38.500 ;
        RECT 116.420 35.850 118.210 37.970 ;
        RECT 118.750 35.860 119.390 38.520 ;
        RECT 119.940 35.850 121.710 37.970 ;
        RECT 122.260 35.860 122.870 38.520 ;
        RECT 123.430 38.510 126.390 39.120 ;
        RECT 126.930 38.520 129.900 39.120 ;
        RECT 130.430 38.790 133.425 39.150 ;
        RECT 130.430 38.520 133.430 38.790 ;
        RECT 123.450 37.965 125.200 37.970 ;
        RECT 123.450 35.860 125.210 37.965 ;
        RECT 125.770 35.860 126.390 38.510 ;
        RECT 126.960 35.860 128.730 37.970 ;
        RECT 129.290 35.860 129.900 38.520 ;
        RECT 130.470 37.960 131.060 37.965 ;
        RECT 131.640 37.960 132.230 37.965 ;
        RECT 130.470 35.860 132.230 37.960 ;
        RECT 132.780 35.860 133.430 38.520 ;
        RECT 133.980 35.860 135.740 37.970 ;
        RECT 136.320 35.580 137.720 48.820 ;
        RECT 105.090 35.120 137.720 35.580 ;
        RECT 20.050 31.700 133.200 33.700 ;
        RECT 20.400 31.500 24.650 31.700 ;
        RECT 20.400 30.900 95.200 31.500 ;
        RECT 20.400 23.400 21.000 30.900 ;
        RECT 21.850 30.570 22.450 30.600 ;
        RECT 25.990 30.570 26.590 30.600 ;
        RECT 35.630 30.570 36.230 30.600 ;
        RECT 45.270 30.570 45.870 30.600 ;
        RECT 54.910 30.570 55.510 30.600 ;
        RECT 64.550 30.570 65.150 30.600 ;
        RECT 74.190 30.570 74.790 30.600 ;
        RECT 81.300 30.570 81.900 30.605 ;
        RECT 21.650 30.340 22.650 30.570 ;
        RECT 23.290 30.340 32.290 30.570 ;
        RECT 32.930 30.340 41.930 30.570 ;
        RECT 42.570 30.340 51.570 30.570 ;
        RECT 52.210 30.340 61.210 30.570 ;
        RECT 61.850 30.340 70.850 30.570 ;
        RECT 71.490 30.340 80.490 30.570 ;
        RECT 81.130 30.340 82.130 30.570 ;
        RECT 21.850 30.310 22.450 30.340 ;
        RECT 25.990 30.310 26.590 30.340 ;
        RECT 35.630 30.310 36.230 30.340 ;
        RECT 45.270 30.310 45.870 30.340 ;
        RECT 54.910 30.310 55.510 30.340 ;
        RECT 64.550 30.310 65.150 30.340 ;
        RECT 74.190 30.310 74.790 30.340 ;
        RECT 81.300 30.310 81.900 30.340 ;
        RECT 21.215 28.900 21.445 30.290 ;
        RECT 21.150 28.400 21.550 28.900 ;
        RECT 21.215 27.330 21.445 28.400 ;
        RECT 22.855 27.330 23.085 30.290 ;
        RECT 32.495 27.330 32.725 30.290 ;
        RECT 42.135 27.330 42.365 30.290 ;
        RECT 51.775 27.330 52.005 30.290 ;
        RECT 61.415 27.330 61.645 30.290 ;
        RECT 71.055 27.330 71.285 30.290 ;
        RECT 80.695 27.330 80.925 30.290 ;
        RECT 82.335 29.100 82.565 30.290 ;
        RECT 82.200 28.600 82.650 29.100 ;
        RECT 82.335 27.330 82.565 28.600 ;
        RECT 82.800 28.500 83.400 30.900 ;
        RECT 84.900 30.585 85.500 30.650 ;
        RECT 84.040 30.355 94.000 30.585 ;
        RECT 84.900 30.350 85.500 30.355 ;
        RECT 83.760 30.100 83.990 30.150 ;
        RECT 94.050 30.100 94.280 30.150 ;
        RECT 83.650 29.200 84.050 30.100 ;
        RECT 94.000 29.200 94.400 30.100 ;
        RECT 83.760 29.150 83.990 29.200 ;
        RECT 94.050 29.150 94.280 29.200 ;
        RECT 84.900 28.945 85.500 28.950 ;
        RECT 84.040 28.715 94.000 28.945 ;
        RECT 84.900 28.650 85.500 28.715 ;
        RECT 94.600 28.500 95.200 30.900 ;
        RECT 82.800 27.900 95.200 28.500 ;
        RECT 96.150 30.900 133.200 31.500 ;
        RECT 21.850 27.280 22.450 27.310 ;
        RECT 28.990 27.280 29.590 27.310 ;
        RECT 38.630 27.280 39.230 27.310 ;
        RECT 48.270 27.280 48.870 27.310 ;
        RECT 57.910 27.280 58.510 27.310 ;
        RECT 67.550 27.280 68.150 27.310 ;
        RECT 77.190 27.280 77.790 27.310 ;
        RECT 81.300 27.280 81.900 27.315 ;
        RECT 21.650 27.050 22.650 27.280 ;
        RECT 23.290 27.050 32.290 27.280 ;
        RECT 32.930 27.050 41.930 27.280 ;
        RECT 42.570 27.050 51.570 27.280 ;
        RECT 52.210 27.050 61.210 27.280 ;
        RECT 61.850 27.050 70.850 27.280 ;
        RECT 71.490 27.050 80.490 27.280 ;
        RECT 81.130 27.050 82.130 27.280 ;
        RECT 21.850 27.020 22.450 27.050 ;
        RECT 28.990 27.020 29.590 27.050 ;
        RECT 38.630 27.020 39.230 27.050 ;
        RECT 48.270 27.020 48.870 27.050 ;
        RECT 57.910 27.020 58.510 27.050 ;
        RECT 67.550 27.020 68.150 27.050 ;
        RECT 77.190 27.020 77.790 27.050 ;
        RECT 81.300 27.020 81.900 27.050 ;
        RECT 21.215 25.800 21.445 27.000 ;
        RECT 21.150 25.300 21.550 25.800 ;
        RECT 21.215 24.040 21.445 25.300 ;
        RECT 22.855 24.040 23.085 27.000 ;
        RECT 32.495 24.040 32.725 27.000 ;
        RECT 42.135 24.040 42.365 27.000 ;
        RECT 51.775 24.040 52.005 27.000 ;
        RECT 61.415 24.040 61.645 27.000 ;
        RECT 71.055 24.040 71.285 27.000 ;
        RECT 80.695 24.040 80.925 27.000 ;
        RECT 82.335 25.800 82.565 27.000 ;
        RECT 82.200 25.300 82.650 25.800 ;
        RECT 82.335 24.040 82.565 25.300 ;
        RECT 21.850 23.990 22.450 24.020 ;
        RECT 25.990 23.990 26.590 24.020 ;
        RECT 35.630 23.990 36.230 24.020 ;
        RECT 45.270 23.990 45.870 24.020 ;
        RECT 54.910 23.990 55.510 24.020 ;
        RECT 64.550 23.990 65.150 24.020 ;
        RECT 74.190 23.990 74.790 24.020 ;
        RECT 81.300 23.990 81.900 24.020 ;
        RECT 21.650 23.760 22.650 23.990 ;
        RECT 23.290 23.760 32.290 23.990 ;
        RECT 32.930 23.760 41.930 23.990 ;
        RECT 42.570 23.760 51.570 23.990 ;
        RECT 52.210 23.760 61.210 23.990 ;
        RECT 61.850 23.760 70.850 23.990 ;
        RECT 71.490 23.760 80.490 23.990 ;
        RECT 81.130 23.760 82.130 23.990 ;
        RECT 21.850 23.730 22.450 23.760 ;
        RECT 25.990 23.730 26.590 23.760 ;
        RECT 35.630 23.730 36.230 23.760 ;
        RECT 45.270 23.730 45.870 23.760 ;
        RECT 54.910 23.730 55.510 23.760 ;
        RECT 64.550 23.730 65.150 23.760 ;
        RECT 74.190 23.730 74.790 23.760 ;
        RECT 81.300 23.725 81.900 23.760 ;
        RECT 82.800 23.400 83.400 27.900 ;
        RECT 96.150 27.000 96.750 30.900 ;
        RECT 97.510 30.350 98.470 30.580 ;
        RECT 100.200 30.490 100.800 30.520 ;
        RECT 102.190 30.490 102.790 30.520 ;
        RECT 105.740 30.490 106.340 30.520 ;
        RECT 109.290 30.490 109.890 30.520 ;
        RECT 112.840 30.490 113.440 30.520 ;
        RECT 115.950 30.490 116.550 30.520 ;
        RECT 99.940 30.260 100.940 30.490 ;
        RECT 101.490 30.260 104.490 30.490 ;
        RECT 105.040 30.260 108.040 30.490 ;
        RECT 108.590 30.260 111.590 30.490 ;
        RECT 112.140 30.260 115.140 30.490 ;
        RECT 115.690 30.260 116.690 30.490 ;
        RECT 100.200 30.230 100.800 30.260 ;
        RECT 102.190 30.230 102.790 30.260 ;
        RECT 105.740 30.230 106.340 30.260 ;
        RECT 109.290 30.230 109.890 30.260 ;
        RECT 112.840 30.230 113.440 30.260 ;
        RECT 115.950 30.230 116.550 30.260 ;
        RECT 97.230 27.450 97.460 30.190 ;
        RECT 98.520 28.300 98.750 30.190 ;
        RECT 99.550 28.900 99.780 30.210 ;
        RECT 99.300 28.400 99.900 28.900 ;
        RECT 20.400 22.800 83.400 23.400 ;
        RECT 84.200 26.400 96.750 27.000 ;
        RECT 97.150 26.950 97.550 27.450 ;
        RECT 98.400 27.150 99.000 28.300 ;
        RECT 99.550 27.250 99.780 28.400 ;
        RECT 101.100 27.250 101.330 30.210 ;
        RECT 104.650 27.250 104.880 30.210 ;
        RECT 108.200 27.250 108.430 30.210 ;
        RECT 111.750 27.250 111.980 30.210 ;
        RECT 115.300 27.250 115.530 30.210 ;
        RECT 116.850 28.950 117.080 30.210 ;
        RECT 117.680 29.020 119.785 30.330 ;
        RECT 129.975 29.020 132.080 30.330 ;
        RECT 116.800 28.450 117.350 28.950 ;
        RECT 116.850 27.250 117.080 28.450 ;
        RECT 100.200 27.200 100.800 27.230 ;
        RECT 103.190 27.200 103.790 27.230 ;
        RECT 106.740 27.200 107.340 27.230 ;
        RECT 110.290 27.200 110.890 27.230 ;
        RECT 113.835 27.200 114.435 27.230 ;
        RECT 115.950 27.200 116.550 27.230 ;
        RECT 84.200 22.750 84.800 26.400 ;
        RECT 86.100 25.990 86.700 26.050 ;
        RECT 85.490 25.760 95.490 25.990 ;
        RECT 86.100 25.750 86.700 25.760 ;
        RECT 85.100 25.600 85.330 25.710 ;
        RECT 84.950 24.900 85.400 25.600 ;
        RECT 85.100 24.750 85.330 24.900 ;
        RECT 95.650 24.750 95.880 25.710 ;
        RECT 97.230 25.190 97.460 26.950 ;
        RECT 98.520 25.190 98.750 27.150 ;
        RECT 99.940 26.970 100.940 27.200 ;
        RECT 101.490 26.970 104.490 27.200 ;
        RECT 105.040 26.970 108.040 27.200 ;
        RECT 108.590 26.970 111.590 27.200 ;
        RECT 112.140 26.970 115.140 27.200 ;
        RECT 115.690 26.970 116.690 27.200 ;
        RECT 117.680 27.130 119.785 28.440 ;
        RECT 129.975 27.130 132.080 28.440 ;
        RECT 100.200 26.940 100.800 26.970 ;
        RECT 103.190 26.940 103.790 26.970 ;
        RECT 106.740 26.940 107.340 26.970 ;
        RECT 110.290 26.940 110.890 26.970 ;
        RECT 113.835 26.940 114.435 26.970 ;
        RECT 115.950 26.940 116.550 26.970 ;
        RECT 99.550 25.650 99.780 26.920 ;
        RECT 99.300 25.150 99.900 25.650 ;
        RECT 97.600 25.030 98.200 25.100 ;
        RECT 97.510 24.800 98.470 25.030 ;
        RECT 93.900 24.700 94.500 24.750 ;
        RECT 85.490 24.470 95.490 24.700 ;
        RECT 97.600 24.600 98.200 24.800 ;
        RECT 93.900 24.450 94.500 24.470 ;
        RECT 85.100 24.300 85.330 24.420 ;
        RECT 84.950 23.600 85.400 24.300 ;
        RECT 85.100 23.460 85.330 23.600 ;
        RECT 95.650 23.460 95.880 24.420 ;
        RECT 99.550 23.960 99.780 25.150 ;
        RECT 101.100 23.960 101.330 26.920 ;
        RECT 104.650 23.960 104.880 26.920 ;
        RECT 108.200 23.960 108.430 26.920 ;
        RECT 111.750 23.960 111.980 26.920 ;
        RECT 115.300 23.960 115.530 26.920 ;
        RECT 116.850 25.700 117.080 26.920 ;
        RECT 116.800 25.200 117.350 25.700 ;
        RECT 117.680 25.240 119.785 26.550 ;
        RECT 129.975 25.240 132.080 26.550 ;
        RECT 116.850 23.960 117.080 25.200 ;
        RECT 100.200 23.910 100.800 23.940 ;
        RECT 102.190 23.910 102.790 23.940 ;
        RECT 105.740 23.910 106.340 23.940 ;
        RECT 109.290 23.910 109.890 23.940 ;
        RECT 112.840 23.910 113.440 23.940 ;
        RECT 115.950 23.910 116.550 23.940 ;
        RECT 99.940 23.680 100.940 23.910 ;
        RECT 101.490 23.680 104.490 23.910 ;
        RECT 105.040 23.680 108.040 23.910 ;
        RECT 108.590 23.680 111.590 23.910 ;
        RECT 112.140 23.680 115.140 23.910 ;
        RECT 115.690 23.680 116.690 23.910 ;
        RECT 100.200 23.650 100.800 23.680 ;
        RECT 102.190 23.650 102.790 23.680 ;
        RECT 105.740 23.650 106.340 23.680 ;
        RECT 109.290 23.650 109.890 23.680 ;
        RECT 112.840 23.650 113.440 23.680 ;
        RECT 115.950 23.650 116.550 23.680 ;
        RECT 86.100 23.410 86.700 23.450 ;
        RECT 85.490 23.180 95.490 23.410 ;
        RECT 117.680 23.350 119.785 24.660 ;
        RECT 129.975 23.350 132.080 24.660 ;
        RECT 86.100 23.150 86.700 23.180 ;
        RECT 132.600 22.750 133.200 30.900 ;
        RECT 84.200 22.150 133.200 22.750 ;
        RECT 84.200 21.950 85.200 22.150 ;
        RECT 20.050 19.950 133.200 21.950 ;
        RECT 22.200 17.650 23.200 19.950 ;
        RECT 20.400 17.050 134.250 17.650 ;
        RECT 20.400 5.600 21.000 17.050 ;
        RECT 21.850 16.580 22.450 16.610 ;
        RECT 27.650 16.580 28.250 16.610 ;
        RECT 43.200 16.580 43.800 16.610 ;
        RECT 58.750 16.580 59.350 16.610 ;
        RECT 74.300 16.580 74.900 16.610 ;
        RECT 89.850 16.580 90.450 16.610 ;
        RECT 105.400 16.580 106.000 16.610 ;
        RECT 120.950 16.580 121.550 16.610 ;
        RECT 132.250 16.580 132.850 16.610 ;
        RECT 21.650 16.350 22.650 16.580 ;
        RECT 23.200 16.350 38.200 16.580 ;
        RECT 38.750 16.350 53.750 16.580 ;
        RECT 54.300 16.350 69.300 16.580 ;
        RECT 69.850 16.350 84.850 16.580 ;
        RECT 85.400 16.350 100.400 16.580 ;
        RECT 100.950 16.350 115.950 16.580 ;
        RECT 116.500 16.350 131.500 16.580 ;
        RECT 132.050 16.350 133.050 16.580 ;
        RECT 21.850 16.320 22.450 16.350 ;
        RECT 27.650 16.320 28.250 16.350 ;
        RECT 43.200 16.320 43.800 16.350 ;
        RECT 58.750 16.320 59.350 16.350 ;
        RECT 74.300 16.320 74.900 16.350 ;
        RECT 89.850 16.320 90.450 16.350 ;
        RECT 105.400 16.320 106.000 16.350 ;
        RECT 120.950 16.320 121.550 16.350 ;
        RECT 132.250 16.320 132.850 16.350 ;
        RECT 21.260 16.150 21.490 16.300 ;
        RECT 21.150 15.450 21.600 16.150 ;
        RECT 21.260 15.340 21.490 15.450 ;
        RECT 22.810 15.340 23.040 16.300 ;
        RECT 38.360 15.340 38.590 16.300 ;
        RECT 53.910 15.340 54.140 16.300 ;
        RECT 69.460 15.340 69.690 16.300 ;
        RECT 85.010 15.340 85.240 16.300 ;
        RECT 100.560 15.340 100.790 16.300 ;
        RECT 116.110 15.340 116.340 16.300 ;
        RECT 131.660 15.340 131.890 16.300 ;
        RECT 133.210 16.150 133.440 16.300 ;
        RECT 133.050 15.450 133.500 16.150 ;
        RECT 133.210 15.340 133.440 15.450 ;
        RECT 21.850 15.290 22.450 15.320 ;
        RECT 32.650 15.290 33.250 15.320 ;
        RECT 48.200 15.290 48.800 15.320 ;
        RECT 63.750 15.290 64.350 15.320 ;
        RECT 79.300 15.290 79.900 15.320 ;
        RECT 94.850 15.290 95.450 15.320 ;
        RECT 110.400 15.290 111.000 15.320 ;
        RECT 125.950 15.290 126.550 15.320 ;
        RECT 132.250 15.290 132.850 15.320 ;
        RECT 21.650 15.060 22.650 15.290 ;
        RECT 23.200 15.060 38.200 15.290 ;
        RECT 38.750 15.060 53.750 15.290 ;
        RECT 54.300 15.060 69.300 15.290 ;
        RECT 69.850 15.060 84.850 15.290 ;
        RECT 85.400 15.060 100.400 15.290 ;
        RECT 100.950 15.060 115.950 15.290 ;
        RECT 116.500 15.060 131.500 15.290 ;
        RECT 132.050 15.060 133.050 15.290 ;
        RECT 21.850 15.030 22.450 15.060 ;
        RECT 32.650 15.030 33.250 15.060 ;
        RECT 48.200 15.030 48.800 15.060 ;
        RECT 63.750 15.030 64.350 15.060 ;
        RECT 79.300 15.030 79.900 15.060 ;
        RECT 94.850 15.030 95.450 15.060 ;
        RECT 110.400 15.030 111.000 15.060 ;
        RECT 125.950 15.030 126.550 15.060 ;
        RECT 132.250 15.030 132.850 15.060 ;
        RECT 21.260 14.900 21.490 15.010 ;
        RECT 21.150 14.200 21.600 14.900 ;
        RECT 21.260 14.050 21.490 14.200 ;
        RECT 22.810 14.050 23.040 15.010 ;
        RECT 38.360 14.050 38.590 15.010 ;
        RECT 53.910 14.050 54.140 15.010 ;
        RECT 69.460 14.050 69.690 15.010 ;
        RECT 85.010 14.050 85.240 15.010 ;
        RECT 100.560 14.050 100.790 15.010 ;
        RECT 116.110 14.050 116.340 15.010 ;
        RECT 131.660 14.050 131.890 15.010 ;
        RECT 133.210 14.900 133.440 15.010 ;
        RECT 133.050 14.200 133.500 14.900 ;
        RECT 133.210 14.050 133.440 14.200 ;
        RECT 21.850 14.000 22.450 14.030 ;
        RECT 27.650 14.000 28.250 14.030 ;
        RECT 43.200 14.000 43.800 14.030 ;
        RECT 58.750 14.000 59.350 14.030 ;
        RECT 74.300 14.000 74.900 14.030 ;
        RECT 89.850 14.000 90.450 14.030 ;
        RECT 105.400 14.000 106.000 14.030 ;
        RECT 120.950 14.000 121.550 14.030 ;
        RECT 132.250 14.000 132.850 14.030 ;
        RECT 21.650 13.770 22.650 14.000 ;
        RECT 23.200 13.770 38.200 14.000 ;
        RECT 38.750 13.770 53.750 14.000 ;
        RECT 54.300 13.770 69.300 14.000 ;
        RECT 69.850 13.770 84.850 14.000 ;
        RECT 85.400 13.770 100.400 14.000 ;
        RECT 100.950 13.770 115.950 14.000 ;
        RECT 116.500 13.770 131.500 14.000 ;
        RECT 132.050 13.770 133.050 14.000 ;
        RECT 21.850 13.740 22.450 13.770 ;
        RECT 27.650 13.740 28.250 13.770 ;
        RECT 43.200 13.740 43.800 13.770 ;
        RECT 58.750 13.740 59.350 13.770 ;
        RECT 74.300 13.740 74.900 13.770 ;
        RECT 89.850 13.740 90.450 13.770 ;
        RECT 105.400 13.740 106.000 13.770 ;
        RECT 120.950 13.740 121.550 13.770 ;
        RECT 132.250 13.740 132.850 13.770 ;
        RECT 21.260 13.600 21.490 13.720 ;
        RECT 21.150 12.900 21.600 13.600 ;
        RECT 21.260 12.760 21.490 12.900 ;
        RECT 22.810 12.760 23.040 13.720 ;
        RECT 38.360 12.760 38.590 13.720 ;
        RECT 53.910 12.760 54.140 13.720 ;
        RECT 69.460 12.760 69.690 13.720 ;
        RECT 85.010 12.760 85.240 13.720 ;
        RECT 100.560 12.760 100.790 13.720 ;
        RECT 116.110 12.760 116.340 13.720 ;
        RECT 131.660 12.760 131.890 13.720 ;
        RECT 133.210 13.600 133.440 13.720 ;
        RECT 133.050 12.900 133.500 13.600 ;
        RECT 133.210 12.760 133.440 12.900 ;
        RECT 21.850 12.710 22.450 12.740 ;
        RECT 32.650 12.710 33.250 12.740 ;
        RECT 48.200 12.710 48.800 12.740 ;
        RECT 63.750 12.710 64.350 12.740 ;
        RECT 79.300 12.710 79.900 12.740 ;
        RECT 94.850 12.710 95.450 12.740 ;
        RECT 110.400 12.710 111.000 12.740 ;
        RECT 125.950 12.710 126.550 12.740 ;
        RECT 132.250 12.710 132.850 12.740 ;
        RECT 21.650 12.480 22.650 12.710 ;
        RECT 23.200 12.480 38.200 12.710 ;
        RECT 38.750 12.480 53.750 12.710 ;
        RECT 54.300 12.480 69.300 12.710 ;
        RECT 69.850 12.480 84.850 12.710 ;
        RECT 85.400 12.480 100.400 12.710 ;
        RECT 100.950 12.480 115.950 12.710 ;
        RECT 116.500 12.480 131.500 12.710 ;
        RECT 132.050 12.480 133.050 12.710 ;
        RECT 21.850 12.450 22.450 12.480 ;
        RECT 32.650 12.450 33.250 12.480 ;
        RECT 48.200 12.450 48.800 12.480 ;
        RECT 63.750 12.450 64.350 12.480 ;
        RECT 79.300 12.450 79.900 12.480 ;
        RECT 94.850 12.450 95.450 12.480 ;
        RECT 110.400 12.450 111.000 12.480 ;
        RECT 125.950 12.450 126.550 12.480 ;
        RECT 132.250 12.450 132.850 12.480 ;
        RECT 21.260 12.300 21.490 12.430 ;
        RECT 21.150 11.600 21.600 12.300 ;
        RECT 21.260 11.470 21.490 11.600 ;
        RECT 22.810 11.470 23.040 12.430 ;
        RECT 38.360 11.470 38.590 12.430 ;
        RECT 53.910 11.470 54.140 12.430 ;
        RECT 69.460 11.470 69.690 12.430 ;
        RECT 85.010 11.470 85.240 12.430 ;
        RECT 100.560 11.470 100.790 12.430 ;
        RECT 116.110 11.470 116.340 12.430 ;
        RECT 131.660 11.470 131.890 12.430 ;
        RECT 133.210 12.300 133.440 12.430 ;
        RECT 133.050 11.600 133.500 12.300 ;
        RECT 133.210 11.470 133.440 11.600 ;
        RECT 21.850 11.420 22.450 11.450 ;
        RECT 27.650 11.420 28.250 11.450 ;
        RECT 43.200 11.420 43.800 11.450 ;
        RECT 58.750 11.420 59.350 11.450 ;
        RECT 74.300 11.420 74.900 11.450 ;
        RECT 89.850 11.420 90.450 11.450 ;
        RECT 105.400 11.420 106.000 11.450 ;
        RECT 120.950 11.420 121.550 11.450 ;
        RECT 132.250 11.420 132.850 11.450 ;
        RECT 21.650 11.190 22.650 11.420 ;
        RECT 23.200 11.190 38.200 11.420 ;
        RECT 38.750 11.190 53.750 11.420 ;
        RECT 54.300 11.190 69.300 11.420 ;
        RECT 69.850 11.190 84.850 11.420 ;
        RECT 85.400 11.190 100.400 11.420 ;
        RECT 100.950 11.190 115.950 11.420 ;
        RECT 116.500 11.190 131.500 11.420 ;
        RECT 132.050 11.190 133.050 11.420 ;
        RECT 21.850 11.160 22.450 11.190 ;
        RECT 27.650 11.160 28.250 11.190 ;
        RECT 43.200 11.160 43.800 11.190 ;
        RECT 58.750 11.160 59.350 11.190 ;
        RECT 74.300 11.160 74.900 11.190 ;
        RECT 89.850 11.160 90.450 11.190 ;
        RECT 105.400 11.160 106.000 11.190 ;
        RECT 120.950 11.160 121.550 11.190 ;
        RECT 132.250 11.160 132.850 11.190 ;
        RECT 21.260 11.000 21.490 11.140 ;
        RECT 21.150 10.300 21.600 11.000 ;
        RECT 21.260 10.180 21.490 10.300 ;
        RECT 22.810 10.180 23.040 11.140 ;
        RECT 38.360 10.180 38.590 11.140 ;
        RECT 53.910 10.180 54.140 11.140 ;
        RECT 69.460 10.180 69.690 11.140 ;
        RECT 85.010 10.180 85.240 11.140 ;
        RECT 100.560 10.180 100.790 11.140 ;
        RECT 116.110 10.180 116.340 11.140 ;
        RECT 131.660 10.180 131.890 11.140 ;
        RECT 133.210 11.050 133.440 11.140 ;
        RECT 133.050 10.350 133.500 11.050 ;
        RECT 133.210 10.180 133.440 10.350 ;
        RECT 21.850 10.130 22.450 10.160 ;
        RECT 32.650 10.130 33.250 10.160 ;
        RECT 48.200 10.130 48.800 10.160 ;
        RECT 63.750 10.130 64.350 10.160 ;
        RECT 79.300 10.130 79.900 10.160 ;
        RECT 94.850 10.130 95.450 10.160 ;
        RECT 110.400 10.130 111.000 10.160 ;
        RECT 125.950 10.130 126.550 10.160 ;
        RECT 132.250 10.130 132.850 10.160 ;
        RECT 21.650 9.900 22.650 10.130 ;
        RECT 23.200 9.900 38.200 10.130 ;
        RECT 38.750 9.900 53.750 10.130 ;
        RECT 54.300 9.900 69.300 10.130 ;
        RECT 69.850 9.900 84.850 10.130 ;
        RECT 85.400 9.900 100.400 10.130 ;
        RECT 100.950 9.900 115.950 10.130 ;
        RECT 116.500 9.900 131.500 10.130 ;
        RECT 132.050 9.900 133.050 10.130 ;
        RECT 21.850 9.870 22.450 9.900 ;
        RECT 32.650 9.870 33.250 9.900 ;
        RECT 48.200 9.870 48.800 9.900 ;
        RECT 63.750 9.870 64.350 9.900 ;
        RECT 79.300 9.870 79.900 9.900 ;
        RECT 94.850 9.870 95.450 9.900 ;
        RECT 110.400 9.870 111.000 9.900 ;
        RECT 125.950 9.870 126.550 9.900 ;
        RECT 132.250 9.870 132.850 9.900 ;
        RECT 21.260 9.700 21.490 9.850 ;
        RECT 21.150 9.000 21.600 9.700 ;
        RECT 21.260 8.890 21.490 9.000 ;
        RECT 22.810 8.890 23.040 9.850 ;
        RECT 38.360 8.890 38.590 9.850 ;
        RECT 53.910 8.890 54.140 9.850 ;
        RECT 69.460 8.890 69.690 9.850 ;
        RECT 85.010 8.890 85.240 9.850 ;
        RECT 100.560 8.890 100.790 9.850 ;
        RECT 116.110 8.890 116.340 9.850 ;
        RECT 131.660 8.890 131.890 9.850 ;
        RECT 133.210 9.750 133.440 9.850 ;
        RECT 133.050 9.050 133.500 9.750 ;
        RECT 133.210 8.890 133.440 9.050 ;
        RECT 21.850 8.840 22.450 8.870 ;
        RECT 27.650 8.840 28.250 8.870 ;
        RECT 43.200 8.840 43.800 8.870 ;
        RECT 58.750 8.840 59.350 8.870 ;
        RECT 74.300 8.840 74.900 8.870 ;
        RECT 89.850 8.840 90.450 8.870 ;
        RECT 105.400 8.840 106.000 8.870 ;
        RECT 120.950 8.840 121.550 8.870 ;
        RECT 132.250 8.840 132.850 8.870 ;
        RECT 21.650 8.610 22.650 8.840 ;
        RECT 23.200 8.610 38.200 8.840 ;
        RECT 38.750 8.610 53.750 8.840 ;
        RECT 54.300 8.610 69.300 8.840 ;
        RECT 69.850 8.610 84.850 8.840 ;
        RECT 85.400 8.610 100.400 8.840 ;
        RECT 100.950 8.610 115.950 8.840 ;
        RECT 116.500 8.610 131.500 8.840 ;
        RECT 132.050 8.610 133.050 8.840 ;
        RECT 21.850 8.580 22.450 8.610 ;
        RECT 27.650 8.580 28.250 8.610 ;
        RECT 43.200 8.580 43.800 8.610 ;
        RECT 58.750 8.580 59.350 8.610 ;
        RECT 74.300 8.580 74.900 8.610 ;
        RECT 89.850 8.580 90.450 8.610 ;
        RECT 105.400 8.580 106.000 8.610 ;
        RECT 120.950 8.580 121.550 8.610 ;
        RECT 132.250 8.580 132.850 8.610 ;
        RECT 21.260 8.450 21.490 8.560 ;
        RECT 21.150 7.750 21.600 8.450 ;
        RECT 21.260 7.600 21.490 7.750 ;
        RECT 22.810 7.600 23.040 8.560 ;
        RECT 38.360 7.600 38.590 8.560 ;
        RECT 53.910 7.600 54.140 8.560 ;
        RECT 69.460 7.600 69.690 8.560 ;
        RECT 85.010 7.600 85.240 8.560 ;
        RECT 100.560 7.600 100.790 8.560 ;
        RECT 116.110 7.600 116.340 8.560 ;
        RECT 131.660 7.600 131.890 8.560 ;
        RECT 133.210 8.450 133.440 8.560 ;
        RECT 133.050 7.750 133.500 8.450 ;
        RECT 133.210 7.600 133.440 7.750 ;
        RECT 21.850 7.550 22.450 7.580 ;
        RECT 32.650 7.550 33.250 7.580 ;
        RECT 48.200 7.550 48.800 7.580 ;
        RECT 63.750 7.550 64.350 7.580 ;
        RECT 79.300 7.550 79.900 7.580 ;
        RECT 94.850 7.550 95.450 7.580 ;
        RECT 110.400 7.550 111.000 7.580 ;
        RECT 125.950 7.550 126.550 7.580 ;
        RECT 132.250 7.550 132.850 7.580 ;
        RECT 21.650 7.320 22.650 7.550 ;
        RECT 23.200 7.320 38.200 7.550 ;
        RECT 38.750 7.320 53.750 7.550 ;
        RECT 54.300 7.320 69.300 7.550 ;
        RECT 69.850 7.320 84.850 7.550 ;
        RECT 85.400 7.320 100.400 7.550 ;
        RECT 100.950 7.320 115.950 7.550 ;
        RECT 116.500 7.320 131.500 7.550 ;
        RECT 132.050 7.320 133.050 7.550 ;
        RECT 21.850 7.290 22.450 7.320 ;
        RECT 32.650 7.290 33.250 7.320 ;
        RECT 48.200 7.290 48.800 7.320 ;
        RECT 63.750 7.290 64.350 7.320 ;
        RECT 79.300 7.290 79.900 7.320 ;
        RECT 94.850 7.290 95.450 7.320 ;
        RECT 110.400 7.290 111.000 7.320 ;
        RECT 125.950 7.290 126.550 7.320 ;
        RECT 132.250 7.290 132.850 7.320 ;
        RECT 21.260 7.150 21.490 7.270 ;
        RECT 21.150 6.450 21.600 7.150 ;
        RECT 21.260 6.310 21.490 6.450 ;
        RECT 22.810 6.310 23.040 7.270 ;
        RECT 38.360 6.310 38.590 7.270 ;
        RECT 53.910 6.310 54.140 7.270 ;
        RECT 69.460 6.310 69.690 7.270 ;
        RECT 85.010 6.310 85.240 7.270 ;
        RECT 100.560 6.310 100.790 7.270 ;
        RECT 116.110 6.310 116.340 7.270 ;
        RECT 131.660 6.310 131.890 7.270 ;
        RECT 133.210 7.150 133.440 7.270 ;
        RECT 133.050 6.450 133.500 7.150 ;
        RECT 133.210 6.310 133.440 6.450 ;
        RECT 21.850 6.260 22.450 6.285 ;
        RECT 27.650 6.260 28.250 6.290 ;
        RECT 43.200 6.260 43.800 6.290 ;
        RECT 58.750 6.260 59.350 6.290 ;
        RECT 74.300 6.260 74.900 6.290 ;
        RECT 89.850 6.260 90.450 6.290 ;
        RECT 105.400 6.260 106.000 6.290 ;
        RECT 120.950 6.260 121.550 6.290 ;
        RECT 132.250 6.260 132.850 6.290 ;
        RECT 21.650 6.030 22.650 6.260 ;
        RECT 23.200 6.030 38.200 6.260 ;
        RECT 38.750 6.030 53.750 6.260 ;
        RECT 54.300 6.030 69.300 6.260 ;
        RECT 69.850 6.030 84.850 6.260 ;
        RECT 85.400 6.030 100.400 6.260 ;
        RECT 100.950 6.030 115.950 6.260 ;
        RECT 116.500 6.030 131.500 6.260 ;
        RECT 132.050 6.030 133.050 6.260 ;
        RECT 21.850 6.000 22.450 6.030 ;
        RECT 27.650 6.000 28.250 6.030 ;
        RECT 43.200 6.000 43.800 6.030 ;
        RECT 58.750 6.000 59.350 6.030 ;
        RECT 74.300 6.000 74.900 6.030 ;
        RECT 89.850 6.000 90.450 6.030 ;
        RECT 105.400 6.000 106.000 6.030 ;
        RECT 120.950 6.000 121.550 6.030 ;
        RECT 132.250 6.000 132.850 6.030 ;
        RECT 133.650 5.600 134.250 17.050 ;
        RECT 20.400 5.000 134.250 5.600 ;
      LAYER met2 ;
        RECT 37.120 158.610 37.400 160.000 ;
        RECT 44.940 158.610 45.220 160.000 ;
        RECT 52.760 158.610 53.040 160.000 ;
        RECT 37.120 158.470 37.790 158.610 ;
        RECT 37.120 158.000 37.400 158.470 ;
        RECT 37.650 154.790 37.790 158.470 ;
        RECT 44.940 158.470 46.070 158.610 ;
        RECT 44.940 158.000 45.220 158.470 ;
        RECT 43.675 155.975 45.215 156.345 ;
        RECT 37.590 154.470 37.850 154.790 ;
        RECT 43.675 150.535 45.215 150.905 ;
        RECT 43.675 145.095 45.215 145.465 ;
        RECT 45.930 141.725 46.070 158.470 ;
        RECT 52.760 158.470 54.810 158.610 ;
        RECT 52.760 158.000 53.040 158.470 ;
        RECT 51.850 153.790 52.110 154.110 ;
        RECT 51.910 146.970 52.050 153.790 ;
        RECT 52.930 153.255 54.470 153.625 ;
        RECT 54.670 153.090 54.810 158.470 ;
        RECT 60.580 158.000 60.860 160.000 ;
        RECT 68.400 158.000 68.680 160.000 ;
        RECT 76.220 158.000 76.500 160.000 ;
        RECT 84.040 158.000 84.320 160.000 ;
        RECT 91.860 158.610 92.140 160.000 ;
        RECT 99.680 158.610 99.960 160.000 ;
        RECT 91.860 158.470 94.370 158.610 ;
        RECT 91.860 158.000 92.140 158.470 ;
        RECT 55.530 153.790 55.790 154.110 ;
        RECT 54.610 152.770 54.870 153.090 ;
        RECT 55.590 152.410 55.730 153.790 ;
        RECT 60.650 153.090 60.790 158.000 ;
        RECT 62.185 155.975 63.725 156.345 ;
        RECT 68.470 153.090 68.610 158.000 ;
        RECT 76.290 155.810 76.430 158.000 ;
        RECT 80.695 155.975 82.235 156.345 ;
        RECT 76.230 155.490 76.490 155.810 ;
        RECT 74.850 154.470 75.110 154.790 ;
        RECT 71.440 153.255 72.980 153.625 ;
        RECT 60.590 152.770 60.850 153.090 ;
        RECT 68.410 152.770 68.670 153.090 ;
        RECT 67.950 152.430 68.210 152.750 ;
        RECT 71.170 152.430 71.430 152.750 ;
        RECT 55.530 152.090 55.790 152.410 ;
        RECT 61.510 152.090 61.770 152.410 ;
        RECT 63.810 152.090 64.070 152.410 ;
        RECT 64.270 152.090 64.530 152.410 ;
        RECT 52.930 147.815 54.470 148.185 ;
        RECT 51.850 146.650 52.110 146.970 ;
        RECT 47.710 146.310 47.970 146.630 ;
        RECT 45.860 141.355 46.140 141.725 ;
        RECT 47.770 141.190 47.910 146.310 ;
        RECT 51.390 145.630 51.650 145.950 ;
        RECT 51.450 141.870 51.590 145.630 ;
        RECT 52.930 142.375 54.470 142.745 ;
        RECT 51.390 141.550 51.650 141.870 ;
        RECT 54.610 141.550 54.870 141.870 ;
        RECT 47.710 140.870 47.970 141.190 ;
        RECT 43.675 139.655 45.215 140.025 ;
        RECT 52.930 136.935 54.470 137.305 ;
        RECT 54.670 136.430 54.810 141.550 ;
        RECT 55.590 138.470 55.730 152.090 ;
        RECT 56.910 151.750 57.170 152.070 ;
        RECT 56.970 149.690 57.110 151.750 ;
        RECT 60.590 151.070 60.850 151.390 ;
        RECT 56.910 149.370 57.170 149.690 ;
        RECT 56.450 145.630 56.710 145.950 ;
        RECT 56.510 144.250 56.650 145.630 ;
        RECT 56.970 144.930 57.110 149.370 ;
        RECT 60.650 149.010 60.790 151.070 ;
        RECT 60.590 148.690 60.850 149.010 ;
        RECT 60.130 148.350 60.390 148.670 ;
        RECT 58.290 146.990 58.550 147.310 ;
        RECT 58.350 146.630 58.490 146.990 ;
        RECT 60.190 146.970 60.330 148.350 ;
        RECT 60.130 146.650 60.390 146.970 ;
        RECT 57.370 146.310 57.630 146.630 ;
        RECT 58.290 146.310 58.550 146.630 ;
        RECT 57.430 144.930 57.570 146.310 ;
        RECT 58.350 145.950 58.490 146.310 ;
        RECT 58.290 145.630 58.550 145.950 ;
        RECT 56.910 144.610 57.170 144.930 ;
        RECT 57.370 144.610 57.630 144.930 ;
        RECT 56.450 143.930 56.710 144.250 ;
        RECT 56.970 142.210 57.110 144.610 ;
        RECT 56.910 141.890 57.170 142.210 ;
        RECT 55.990 141.550 56.250 141.870 ;
        RECT 56.050 139.490 56.190 141.550 ;
        RECT 55.990 139.170 56.250 139.490 ;
        RECT 60.190 138.470 60.330 146.650 ;
        RECT 61.570 146.630 61.710 152.090 ;
        RECT 62.185 150.535 63.725 150.905 ;
        RECT 63.350 148.690 63.610 149.010 ;
        RECT 63.410 147.650 63.550 148.690 ;
        RECT 63.350 147.330 63.610 147.650 ;
        RECT 61.050 146.310 61.310 146.630 ;
        RECT 61.510 146.310 61.770 146.630 ;
        RECT 60.590 143.930 60.850 144.250 ;
        RECT 60.650 138.470 60.790 143.930 ;
        RECT 61.110 141.870 61.250 146.310 ;
        RECT 61.570 142.210 61.710 146.310 ;
        RECT 62.185 145.095 63.725 145.465 ;
        RECT 62.890 144.610 63.150 144.930 ;
        RECT 62.950 143.230 63.090 144.610 ;
        RECT 62.890 142.910 63.150 143.230 ;
        RECT 61.510 141.890 61.770 142.210 ;
        RECT 61.050 141.550 61.310 141.870 ;
        RECT 62.950 141.530 63.090 142.910 ;
        RECT 61.510 141.210 61.770 141.530 ;
        RECT 62.890 141.210 63.150 141.530 ;
        RECT 61.570 139.150 61.710 141.210 ;
        RECT 62.185 139.655 63.725 140.025 ;
        RECT 61.510 138.830 61.770 139.150 ;
        RECT 55.530 138.150 55.790 138.470 ;
        RECT 60.130 138.150 60.390 138.470 ;
        RECT 60.590 138.150 60.850 138.470 ;
        RECT 59.210 137.470 59.470 137.790 ;
        RECT 53.230 136.110 53.490 136.430 ;
        RECT 54.610 136.110 54.870 136.430 ;
        RECT 43.675 134.215 45.215 134.585 ;
        RECT 53.290 133.370 53.430 136.110 ;
        RECT 59.270 135.750 59.410 137.470 ;
        RECT 63.870 136.770 64.010 152.090 ;
        RECT 64.330 150.370 64.470 152.090 ;
        RECT 67.490 151.750 67.750 152.070 ;
        RECT 64.270 150.050 64.530 150.370 ;
        RECT 65.190 149.710 65.450 150.030 ;
        RECT 65.250 147.050 65.390 149.710 ;
        RECT 67.030 148.350 67.290 148.670 ;
        RECT 64.790 146.910 65.390 147.050 ;
        RECT 67.090 147.050 67.230 148.350 ;
        RECT 67.550 147.650 67.690 151.750 ;
        RECT 68.010 150.370 68.150 152.430 ;
        RECT 71.230 150.370 71.370 152.430 ;
        RECT 73.470 151.410 73.730 151.730 ;
        RECT 67.950 150.050 68.210 150.370 ;
        RECT 71.170 150.050 71.430 150.370 ;
        RECT 68.010 147.730 68.150 150.050 ;
        RECT 73.530 150.030 73.670 151.410 ;
        RECT 74.910 151.390 75.050 154.470 ;
        RECT 77.610 151.750 77.870 152.070 ;
        RECT 74.850 151.070 75.110 151.390 ;
        RECT 73.470 149.710 73.730 150.030 ;
        RECT 74.910 149.690 75.050 151.070 ;
        RECT 74.850 149.370 75.110 149.690 ;
        RECT 73.470 149.030 73.730 149.350 ;
        RECT 70.710 148.350 70.970 148.670 ;
        RECT 67.490 147.330 67.750 147.650 ;
        RECT 68.010 147.590 69.070 147.730 ;
        RECT 67.090 146.970 68.610 147.050 ;
        RECT 64.790 146.290 64.930 146.910 ;
        RECT 66.110 146.650 66.370 146.970 ;
        RECT 67.090 146.910 68.670 146.970 ;
        RECT 64.730 145.970 64.990 146.290 ;
        RECT 65.190 145.970 65.450 146.290 ;
        RECT 64.730 143.250 64.990 143.570 ;
        RECT 64.790 142.405 64.930 143.250 ;
        RECT 64.720 142.035 65.000 142.405 ;
        RECT 65.250 141.870 65.390 145.970 ;
        RECT 65.650 145.630 65.910 145.950 ;
        RECT 65.190 141.550 65.450 141.870 ;
        RECT 65.710 141.530 65.850 145.630 ;
        RECT 66.170 142.210 66.310 146.650 ;
        RECT 67.090 145.950 67.230 146.910 ;
        RECT 68.410 146.650 68.670 146.910 ;
        RECT 67.490 146.310 67.750 146.630 ;
        RECT 67.030 145.630 67.290 145.950 ;
        RECT 67.550 144.930 67.690 146.310 ;
        RECT 67.490 144.610 67.750 144.930 ;
        RECT 66.110 141.890 66.370 142.210 ;
        RECT 65.650 141.210 65.910 141.530 ;
        RECT 67.030 141.210 67.290 141.530 ;
        RECT 65.190 140.870 65.450 141.190 ;
        RECT 64.270 140.530 64.530 140.850 ;
        RECT 64.330 139.150 64.470 140.530 ;
        RECT 64.270 138.830 64.530 139.150 ;
        RECT 64.330 138.470 64.470 138.830 ;
        RECT 65.250 138.470 65.390 140.870 ;
        RECT 64.270 138.150 64.530 138.470 ;
        RECT 65.190 138.150 65.450 138.470 ;
        RECT 65.650 138.150 65.910 138.470 ;
        RECT 66.570 138.150 66.830 138.470 ;
        RECT 63.810 136.450 64.070 136.770 ;
        RECT 59.210 135.430 59.470 135.750 ;
        RECT 62.185 134.215 63.725 134.585 ;
        RECT 53.230 133.050 53.490 133.370 ;
        RECT 63.810 132.710 64.070 133.030 ;
        RECT 52.930 131.495 54.470 131.865 ;
        RECT 63.870 131.330 64.010 132.710 ;
        RECT 63.810 131.010 64.070 131.330 ;
        RECT 43.675 128.775 45.215 129.145 ;
        RECT 62.185 128.775 63.725 129.145 ;
        RECT 65.710 127.590 65.850 138.150 ;
        RECT 66.630 136.770 66.770 138.150 ;
        RECT 67.090 137.790 67.230 141.210 ;
        RECT 67.030 137.470 67.290 137.790 ;
        RECT 66.570 136.450 66.830 136.770 ;
        RECT 68.930 136.090 69.070 147.590 ;
        RECT 70.770 146.970 70.910 148.350 ;
        RECT 71.440 147.815 72.980 148.185 ;
        RECT 70.710 146.650 70.970 146.970 ;
        RECT 70.250 146.310 70.510 146.630 ;
        RECT 69.790 145.970 70.050 146.290 ;
        RECT 69.850 144.590 69.990 145.970 ;
        RECT 69.790 144.270 70.050 144.590 ;
        RECT 70.310 141.190 70.450 146.310 ;
        RECT 73.530 145.950 73.670 149.030 ;
        RECT 74.850 148.350 75.110 148.670 ;
        RECT 74.390 146.310 74.650 146.630 ;
        RECT 70.710 145.630 70.970 145.950 ;
        RECT 73.470 145.630 73.730 145.950 ;
        RECT 70.770 142.210 70.910 145.630 ;
        RECT 74.450 143.910 74.590 146.310 ;
        RECT 74.910 144.590 75.050 148.350 ;
        RECT 77.670 147.650 77.810 151.750 ;
        RECT 80.695 150.535 82.235 150.905 ;
        RECT 84.110 150.370 84.250 158.000 ;
        RECT 89.950 153.255 91.490 153.625 ;
        RECT 91.410 152.430 91.670 152.750 ;
        RECT 86.350 152.090 86.610 152.410 ;
        RECT 87.270 152.090 87.530 152.410 ;
        RECT 84.970 151.070 85.230 151.390 ;
        RECT 84.050 150.050 84.310 150.370 ;
        RECT 78.530 148.690 78.790 149.010 ;
        RECT 81.750 148.690 82.010 149.010 ;
        RECT 77.610 147.330 77.870 147.650 ;
        RECT 75.310 146.650 75.570 146.970 ;
        RECT 78.070 146.880 78.330 146.970 ;
        RECT 78.590 146.880 78.730 148.690 ;
        RECT 78.070 146.740 78.730 146.880 ;
        RECT 78.070 146.650 78.330 146.740 ;
        RECT 74.850 144.270 75.110 144.590 ;
        RECT 74.390 143.590 74.650 143.910 ;
        RECT 73.470 143.250 73.730 143.570 ;
        RECT 71.440 142.375 72.980 142.745 ;
        RECT 73.530 142.290 73.670 143.250 ;
        RECT 70.710 141.890 70.970 142.210 ;
        RECT 73.530 142.150 74.130 142.290 ;
        RECT 73.470 141.210 73.730 141.530 ;
        RECT 70.250 140.870 70.510 141.190 ;
        RECT 70.310 139.490 70.450 140.870 ;
        RECT 73.530 140.510 73.670 141.210 ;
        RECT 73.470 140.190 73.730 140.510 ;
        RECT 73.990 139.490 74.130 142.150 ;
        RECT 74.450 140.510 74.590 143.590 ;
        RECT 74.910 142.210 75.050 144.270 ;
        RECT 75.370 143.910 75.510 146.650 ;
        RECT 78.590 145.950 78.730 146.740 ;
        RECT 78.990 146.310 79.250 146.630 ;
        RECT 78.530 145.630 78.790 145.950 ;
        RECT 76.230 144.610 76.490 144.930 ;
        RECT 75.310 143.590 75.570 143.910 ;
        RECT 76.290 142.210 76.430 144.610 ;
        RECT 77.150 143.590 77.410 143.910 ;
        RECT 74.850 141.890 75.110 142.210 ;
        RECT 76.230 141.890 76.490 142.210 ;
        RECT 74.390 140.190 74.650 140.510 ;
        RECT 70.250 139.170 70.510 139.490 ;
        RECT 73.930 139.170 74.190 139.490 ;
        RECT 70.710 138.150 70.970 138.470 ;
        RECT 69.330 137.470 69.590 137.790 ;
        RECT 67.490 135.770 67.750 136.090 ;
        RECT 68.870 135.770 69.130 136.090 ;
        RECT 67.030 135.090 67.290 135.410 ;
        RECT 67.090 132.690 67.230 135.090 ;
        RECT 67.550 133.030 67.690 135.770 ;
        RECT 69.390 135.750 69.530 137.470 ;
        RECT 69.330 135.430 69.590 135.750 ;
        RECT 67.490 132.710 67.750 133.030 ;
        RECT 67.030 132.370 67.290 132.690 ;
        RECT 67.030 129.990 67.290 130.310 ;
        RECT 67.090 128.270 67.230 129.990 ;
        RECT 69.390 129.630 69.530 135.430 ;
        RECT 70.770 133.370 70.910 138.150 ;
        RECT 71.440 136.935 72.980 137.305 ;
        RECT 74.910 135.750 75.050 141.890 ;
        RECT 75.310 141.550 75.570 141.870 ;
        RECT 75.370 136.090 75.510 141.550 ;
        RECT 77.210 141.530 77.350 143.590 ;
        RECT 77.150 141.210 77.410 141.530 ;
        RECT 78.590 140.930 78.730 145.630 ;
        RECT 79.050 141.870 79.190 146.310 ;
        RECT 81.810 146.290 81.950 148.690 ;
        RECT 83.130 147.330 83.390 147.650 ;
        RECT 83.190 146.970 83.330 147.330 ;
        RECT 82.210 146.650 82.470 146.970 ;
        RECT 82.670 146.650 82.930 146.970 ;
        RECT 83.130 146.650 83.390 146.970 ;
        RECT 81.750 145.970 82.010 146.290 ;
        RECT 82.270 145.950 82.410 146.650 ;
        RECT 82.210 145.630 82.470 145.950 ;
        RECT 80.695 145.095 82.235 145.465 ;
        RECT 82.730 144.330 82.870 146.650 ;
        RECT 81.810 144.190 82.870 144.330 ;
        RECT 81.810 143.910 81.950 144.190 ;
        RECT 80.830 143.590 81.090 143.910 ;
        RECT 81.750 143.590 82.010 143.910 ;
        RECT 78.990 141.550 79.250 141.870 ;
        RECT 80.890 141.530 81.030 143.590 ;
        RECT 83.190 143.570 83.330 146.650 ;
        RECT 84.110 146.630 84.250 150.050 ;
        RECT 85.030 149.350 85.170 151.070 ;
        RECT 85.890 149.710 86.150 150.030 ;
        RECT 84.970 149.030 85.230 149.350 ;
        RECT 85.950 146.970 86.090 149.710 ;
        RECT 86.410 149.350 86.550 152.090 ;
        RECT 86.350 149.030 86.610 149.350 ;
        RECT 85.890 146.650 86.150 146.970 ;
        RECT 86.350 146.650 86.610 146.970 ;
        RECT 84.050 146.310 84.310 146.630 ;
        RECT 85.950 145.950 86.090 146.650 ;
        RECT 83.590 145.630 83.850 145.950 ;
        RECT 85.890 145.630 86.150 145.950 ;
        RECT 83.130 143.250 83.390 143.570 ;
        RECT 80.830 141.210 81.090 141.530 ;
        RECT 78.590 140.790 79.190 140.930 ;
        RECT 82.670 140.870 82.930 141.190 ;
        RECT 79.050 140.510 79.190 140.790 ;
        RECT 78.990 140.190 79.250 140.510 ;
        RECT 78.070 137.470 78.330 137.790 ;
        RECT 77.610 136.450 77.870 136.770 ;
        RECT 75.770 136.110 76.030 136.430 ;
        RECT 75.310 135.770 75.570 136.090 ;
        RECT 74.850 135.430 75.110 135.750 ;
        RECT 70.710 133.050 70.970 133.370 ;
        RECT 73.470 132.030 73.730 132.350 ;
        RECT 74.390 132.030 74.650 132.350 ;
        RECT 71.440 131.495 72.980 131.865 ;
        RECT 73.530 130.990 73.670 132.030 ;
        RECT 73.470 130.670 73.730 130.990 ;
        RECT 69.330 129.310 69.590 129.630 ;
        RECT 67.030 127.950 67.290 128.270 ;
        RECT 69.390 127.590 69.530 129.310 ;
        RECT 74.450 127.930 74.590 132.030 ;
        RECT 74.390 127.610 74.650 127.930 ;
        RECT 65.650 127.270 65.910 127.590 ;
        RECT 69.330 127.270 69.590 127.590 ;
        RECT 52.930 126.055 54.470 126.425 ;
        RECT 71.440 126.055 72.980 126.425 ;
        RECT 43.675 123.335 45.215 123.705 ;
        RECT 62.185 123.335 63.725 123.705 ;
        RECT 52.930 120.615 54.470 120.985 ;
        RECT 71.440 120.615 72.980 120.985 ;
        RECT 43.675 117.895 45.215 118.265 ;
        RECT 62.185 117.895 63.725 118.265 ;
        RECT 52.930 115.175 54.470 115.545 ;
        RECT 71.440 115.175 72.980 115.545 ;
        RECT 43.675 112.455 45.215 112.825 ;
        RECT 62.185 112.455 63.725 112.825 ;
        RECT 52.930 109.735 54.470 110.105 ;
        RECT 71.440 109.735 72.980 110.105 ;
        RECT 43.675 107.015 45.215 107.385 ;
        RECT 62.185 107.015 63.725 107.385 ;
        RECT 52.930 104.295 54.470 104.665 ;
        RECT 71.440 104.295 72.980 104.665 ;
        RECT 43.675 101.575 45.215 101.945 ;
        RECT 62.185 101.575 63.725 101.945 ;
        RECT 52.930 98.855 54.470 99.225 ;
        RECT 71.440 98.855 72.980 99.225 ;
        RECT 43.675 96.135 45.215 96.505 ;
        RECT 62.185 96.135 63.725 96.505 ;
        RECT 75.830 93.870 75.970 136.110 ;
        RECT 77.670 136.090 77.810 136.450 ;
        RECT 78.130 136.090 78.270 137.470 ;
        RECT 79.050 136.430 79.190 140.190 ;
        RECT 80.695 139.655 82.235 140.025 ;
        RECT 82.730 139.490 82.870 140.870 ;
        RECT 82.670 139.170 82.930 139.490 ;
        RECT 79.450 137.810 79.710 138.130 ;
        RECT 82.210 137.810 82.470 138.130 ;
        RECT 78.990 136.110 79.250 136.430 ;
        RECT 77.610 135.770 77.870 136.090 ;
        RECT 78.070 135.770 78.330 136.090 ;
        RECT 79.510 135.070 79.650 137.810 ;
        RECT 81.750 136.110 82.010 136.430 ;
        RECT 79.910 135.770 80.170 136.090 ;
        RECT 76.230 134.750 76.490 135.070 ;
        RECT 78.530 134.750 78.790 135.070 ;
        RECT 79.450 134.750 79.710 135.070 ;
        RECT 76.290 130.650 76.430 134.750 ;
        RECT 78.590 133.030 78.730 134.750 ;
        RECT 79.970 134.050 80.110 135.770 ;
        RECT 81.810 135.070 81.950 136.110 ;
        RECT 82.270 136.090 82.410 137.810 ;
        RECT 83.190 136.170 83.330 143.250 ;
        RECT 83.650 139.150 83.790 145.630 ;
        RECT 86.410 144.930 86.550 146.650 ;
        RECT 84.510 144.610 84.770 144.930 ;
        RECT 86.350 144.610 86.610 144.930 ;
        RECT 84.570 141.870 84.710 144.610 ;
        RECT 84.510 141.550 84.770 141.870 ;
        RECT 84.050 141.210 84.310 141.530 ;
        RECT 84.970 141.210 85.230 141.530 ;
        RECT 83.590 138.830 83.850 139.150 ;
        RECT 83.190 136.090 83.790 136.170 ;
        RECT 82.210 135.770 82.470 136.090 ;
        RECT 83.190 136.030 83.850 136.090 ;
        RECT 83.590 135.770 83.850 136.030 ;
        RECT 82.670 135.430 82.930 135.750 ;
        RECT 81.750 134.750 82.010 135.070 ;
        RECT 80.695 134.215 82.235 134.585 ;
        RECT 82.730 134.050 82.870 135.430 ;
        RECT 84.110 134.050 84.250 141.210 ;
        RECT 85.030 140.850 85.170 141.210 ;
        RECT 87.330 141.190 87.470 152.090 ;
        RECT 88.650 151.750 88.910 152.070 ;
        RECT 88.710 147.650 88.850 151.750 ;
        RECT 91.470 150.370 91.610 152.430 ;
        RECT 94.230 151.390 94.370 158.470 ;
        RECT 97.910 158.470 99.960 158.610 ;
        RECT 94.170 151.070 94.430 151.390 ;
        RECT 91.410 150.050 91.670 150.370 ;
        RECT 94.230 149.690 94.370 151.070 ;
        RECT 94.170 149.370 94.430 149.690 ;
        RECT 89.110 148.350 89.370 148.670 ;
        RECT 88.650 147.330 88.910 147.650 ;
        RECT 89.170 146.970 89.310 148.350 ;
        RECT 89.950 147.815 91.490 148.185 ;
        RECT 89.110 146.650 89.370 146.970 ;
        RECT 97.910 144.930 98.050 158.470 ;
        RECT 99.680 158.000 99.960 158.470 ;
        RECT 107.500 158.000 107.780 160.000 ;
        RECT 99.205 155.975 100.745 156.345 ;
        RECT 99.205 150.535 100.745 150.905 ;
        RECT 99.205 145.095 100.745 145.465 ;
        RECT 97.850 144.610 98.110 144.930 ;
        RECT 96.010 143.590 96.270 143.910 ;
        RECT 89.950 142.375 91.490 142.745 ;
        RECT 96.070 142.210 96.210 143.590 ;
        RECT 96.010 141.890 96.270 142.210 ;
        RECT 95.550 141.210 95.810 141.530 ;
        RECT 87.270 140.870 87.530 141.190 ;
        RECT 84.970 140.530 85.230 140.850 ;
        RECT 85.030 137.790 85.170 140.530 ;
        RECT 87.330 137.790 87.470 140.870 ;
        RECT 95.610 139.490 95.750 141.210 ;
        RECT 95.550 139.170 95.810 139.490 ;
        RECT 97.910 138.810 98.050 144.610 ;
        RECT 99.205 139.655 100.745 140.025 ;
        RECT 107.570 139.490 107.710 158.000 ;
        RECT 108.460 153.255 110.000 153.625 ;
        RECT 108.460 147.815 110.000 148.185 ;
        RECT 108.460 142.375 110.000 142.745 ;
        RECT 107.510 139.170 107.770 139.490 ;
        RECT 97.850 138.490 98.110 138.810 ;
        RECT 93.250 138.150 93.510 138.470 ;
        RECT 95.090 138.150 95.350 138.470 ;
        RECT 96.010 138.150 96.270 138.470 ;
        RECT 84.970 137.470 85.230 137.790 ;
        RECT 87.270 137.470 87.530 137.790 ;
        RECT 85.030 136.090 85.170 137.470 ;
        RECT 84.970 135.770 85.230 136.090 ;
        RECT 87.330 135.750 87.470 137.470 ;
        RECT 89.950 136.935 91.490 137.305 ;
        RECT 93.310 136.770 93.450 138.150 ;
        RECT 93.250 136.450 93.510 136.770 ;
        RECT 90.030 136.110 90.290 136.430 ;
        RECT 87.270 135.430 87.530 135.750 ;
        RECT 79.910 133.730 80.170 134.050 ;
        RECT 82.670 133.730 82.930 134.050 ;
        RECT 84.050 133.730 84.310 134.050 ;
        RECT 87.330 133.370 87.470 135.430 ;
        RECT 90.090 134.050 90.230 136.110 ;
        RECT 90.030 133.730 90.290 134.050 ;
        RECT 87.270 133.050 87.530 133.370 ;
        RECT 95.150 133.030 95.290 138.150 ;
        RECT 96.070 136.770 96.210 138.150 ;
        RECT 108.460 136.935 110.000 137.305 ;
        RECT 96.010 136.450 96.270 136.770 ;
        RECT 99.205 134.215 100.745 134.585 ;
        RECT 78.070 132.710 78.330 133.030 ;
        RECT 78.530 132.710 78.790 133.030 ;
        RECT 84.050 132.710 84.310 133.030 ;
        RECT 95.090 132.710 95.350 133.030 ;
        RECT 78.130 130.650 78.270 132.710 ;
        RECT 83.590 132.370 83.850 132.690 ;
        RECT 83.650 131.330 83.790 132.370 ;
        RECT 84.110 132.350 84.250 132.710 ;
        RECT 84.050 132.030 84.310 132.350 ;
        RECT 83.590 131.010 83.850 131.330 ;
        RECT 84.110 130.650 84.250 132.030 ;
        RECT 89.950 131.495 91.490 131.865 ;
        RECT 108.460 131.495 110.000 131.865 ;
        RECT 76.230 130.330 76.490 130.650 ;
        RECT 78.070 130.330 78.330 130.650 ;
        RECT 84.050 130.330 84.310 130.650 ;
        RECT 80.695 128.775 82.235 129.145 ;
        RECT 99.205 128.775 100.745 129.145 ;
        RECT 89.950 126.055 91.490 126.425 ;
        RECT 108.460 126.055 110.000 126.425 ;
        RECT 80.695 123.335 82.235 123.705 ;
        RECT 99.205 123.335 100.745 123.705 ;
        RECT 89.950 120.615 91.490 120.985 ;
        RECT 108.460 120.615 110.000 120.985 ;
        RECT 80.695 117.895 82.235 118.265 ;
        RECT 99.205 117.895 100.745 118.265 ;
        RECT 89.950 115.175 91.490 115.545 ;
        RECT 108.460 115.175 110.000 115.545 ;
        RECT 80.695 112.455 82.235 112.825 ;
        RECT 99.205 112.455 100.745 112.825 ;
        RECT 89.950 109.735 91.490 110.105 ;
        RECT 108.460 109.735 110.000 110.105 ;
        RECT 80.695 107.015 82.235 107.385 ;
        RECT 99.205 107.015 100.745 107.385 ;
        RECT 89.950 104.295 91.490 104.665 ;
        RECT 108.460 104.295 110.000 104.665 ;
        RECT 80.695 101.575 82.235 101.945 ;
        RECT 99.205 101.575 100.745 101.945 ;
        RECT 89.950 98.855 91.490 99.225 ;
        RECT 108.460 98.855 110.000 99.225 ;
        RECT 80.695 96.135 82.235 96.505 ;
        RECT 99.205 96.135 100.745 96.505 ;
        RECT 52.930 93.415 54.470 93.785 ;
        RECT 71.440 93.415 72.980 93.785 ;
        RECT 75.370 93.730 75.970 93.870 ;
        RECT 43.675 90.695 45.215 91.065 ;
        RECT 62.185 90.695 63.725 91.065 ;
        RECT 52.930 87.975 54.470 88.345 ;
        RECT 71.440 87.975 72.980 88.345 ;
        RECT 43.675 85.255 45.215 85.625 ;
        RECT 62.185 85.255 63.725 85.625 ;
        RECT 75.370 85.090 75.510 93.730 ;
        RECT 89.950 93.415 91.490 93.785 ;
        RECT 108.460 93.415 110.000 93.785 ;
        RECT 80.695 90.695 82.235 91.065 ;
        RECT 99.205 90.695 100.745 91.065 ;
        RECT 89.950 87.975 91.490 88.345 ;
        RECT 108.460 87.975 110.000 88.345 ;
        RECT 80.695 85.255 82.235 85.625 ;
        RECT 99.205 85.255 100.745 85.625 ;
        RECT 75.310 84.770 75.570 85.090 ;
        RECT 74.850 83.410 75.110 83.730 ;
        RECT 52.930 82.535 54.470 82.905 ;
        RECT 71.440 82.535 72.980 82.905 ;
        RECT 74.910 82.370 75.050 83.410 ;
        RECT 89.950 82.535 91.490 82.905 ;
        RECT 108.460 82.535 110.000 82.905 ;
        RECT 72.550 82.280 72.810 82.370 ;
        RECT 72.150 82.140 72.810 82.280 ;
        RECT 72.150 82.000 72.290 82.140 ;
        RECT 72.550 82.050 72.810 82.140 ;
        RECT 74.850 82.050 75.110 82.370 ;
        RECT 72.080 80.000 72.360 82.000 ;
        RECT 105.000 77.160 107.810 79.050 ;
        RECT 108.990 78.120 109.410 79.010 ;
        RECT 20.550 75.850 23.550 75.955 ;
        RECT 20.550 75.560 23.600 75.850 ;
        RECT 28.750 75.560 29.350 75.850 ;
        RECT 20.550 75.455 23.550 75.560 ;
        RECT 23.870 75.060 24.270 75.560 ;
        RECT 24.800 75.060 26.285 75.560 ;
        RECT 22.750 74.770 23.350 75.060 ;
        RECT 29.750 74.770 30.850 75.060 ;
        RECT 23.750 73.600 25.400 74.100 ;
        RECT 22.750 72.430 23.350 72.720 ;
        RECT 28.750 72.430 29.350 72.720 ;
        RECT 21.750 71.930 23.230 72.035 ;
        RECT 23.850 71.930 24.250 72.430 ;
        RECT 25.900 71.930 26.300 72.430 ;
        RECT 21.750 71.640 23.280 71.930 ;
        RECT 21.750 71.535 23.230 71.640 ;
        RECT 23.850 71.140 24.250 71.640 ;
        RECT 25.900 71.140 26.300 71.640 ;
        RECT 29.750 71.635 30.850 71.930 ;
        RECT 22.680 70.850 23.280 71.140 ;
        RECT 28.750 70.850 29.350 71.140 ;
        RECT 21.750 70.000 23.300 70.500 ;
        RECT 23.850 70.350 24.250 70.850 ;
        RECT 25.900 70.350 26.300 70.850 ;
        RECT 29.750 70.060 30.850 70.350 ;
        RECT 20.300 68.850 21.400 69.850 ;
        RECT 22.750 69.350 26.400 69.850 ;
        RECT 21.750 68.350 39.050 68.850 ;
        RECT 47.730 59.950 48.230 71.500 ;
        RECT 48.550 59.950 49.050 72.900 ;
        RECT 53.190 59.950 53.690 72.900 ;
        RECT 47.600 42.900 48.100 59.000 ;
        RECT 55.440 58.400 55.940 70.920 ;
        RECT 60.080 60.470 60.580 72.950 ;
        RECT 60.075 60.080 60.580 60.470 ;
        RECT 60.080 59.950 60.580 60.080 ;
        RECT 62.330 60.000 62.830 70.920 ;
        RECT 62.330 59.400 62.835 60.000 ;
        RECT 66.970 59.950 67.470 72.950 ;
        RECT 69.220 59.950 69.720 71.500 ;
        RECT 73.860 68.210 74.360 72.950 ;
        RECT 73.855 67.820 74.360 68.210 ;
        RECT 73.860 59.950 74.360 67.820 ;
        RECT 76.110 59.400 76.610 70.920 ;
        RECT 80.750 59.950 81.250 72.950 ;
        RECT 83.000 58.400 83.500 70.920 ;
        RECT 87.640 59.950 88.140 72.950 ;
        RECT 88.460 59.950 88.960 71.500 ;
        RECT 97.750 59.400 98.250 70.500 ;
        RECT 98.750 63.780 99.250 69.930 ;
        RECT 100.150 68.870 100.650 72.900 ;
        RECT 100.450 63.780 100.950 68.470 ;
        RECT 98.700 63.390 99.300 63.780 ;
        RECT 100.400 63.390 101.000 63.780 ;
        RECT 99.540 59.400 99.830 60.000 ;
        RECT 102.120 59.400 102.410 60.000 ;
        RECT 43.950 37.450 44.450 41.950 ;
        RECT 53.850 41.350 54.350 56.250 ;
        RECT 45.725 39.980 46.230 40.370 ;
        RECT 52.275 39.980 52.780 40.370 ;
        RECT 45.725 39.080 46.225 39.980 ;
        RECT 45.725 38.690 46.230 39.080 ;
        RECT 45.725 37.790 46.225 38.690 ;
        RECT 52.275 37.790 52.775 39.980 ;
        RECT 45.725 37.400 46.230 37.790 ;
        RECT 45.725 36.050 46.225 37.400 ;
        RECT 45.725 35.150 46.230 36.050 ;
        RECT 52.275 35.150 52.780 37.790 ;
        RECT 55.275 37.400 55.775 42.950 ;
        RECT 60.100 42.350 60.600 56.300 ;
        RECT 67.600 42.900 68.100 57.000 ;
        RECT 68.600 42.900 69.100 58.000 ;
        RECT 61.825 39.980 62.330 40.370 ;
        RECT 61.825 37.790 62.325 39.980 ;
        RECT 61.825 35.150 62.330 37.790 ;
        RECT 64.825 37.400 65.325 41.950 ;
        RECT 71.375 39.980 71.880 40.370 ;
        RECT 71.375 37.790 71.875 39.980 ;
        RECT 74.375 39.080 74.875 41.950 ;
        RECT 76.100 41.350 76.600 56.300 ;
        RECT 82.350 42.350 82.850 56.300 ;
        RECT 88.600 43.020 89.100 59.000 ;
        RECT 103.550 49.300 104.050 62.850 ;
        RECT 98.250 48.700 98.540 49.300 ;
        RECT 100.830 48.700 101.120 49.300 ;
        RECT 103.410 48.700 104.050 49.300 ;
        RECT 105.080 48.770 107.810 50.070 ;
        RECT 108.140 50.020 108.430 76.850 ;
        RECT 108.995 59.270 109.410 78.120 ;
        RECT 108.610 58.770 109.410 59.270 ;
        RECT 109.720 50.020 110.010 76.840 ;
        RECT 108.140 49.020 110.010 50.020 ;
        RECT 111.840 50.030 112.130 76.860 ;
        RECT 112.580 59.270 112.980 79.010 ;
        RECT 112.320 58.770 112.980 59.270 ;
        RECT 113.420 50.030 113.710 76.850 ;
        RECT 111.840 49.030 113.710 50.030 ;
        RECT 115.550 50.030 115.840 76.860 ;
        RECT 116.310 59.270 116.710 79.010 ;
        RECT 116.020 58.770 116.710 59.270 ;
        RECT 117.130 50.030 117.420 76.850 ;
        RECT 115.550 49.030 117.420 50.030 ;
        RECT 119.260 50.030 119.550 76.860 ;
        RECT 120.020 59.270 120.420 79.010 ;
        RECT 119.730 58.770 120.420 59.270 ;
        RECT 120.840 50.030 121.130 76.850 ;
        RECT 119.260 49.030 121.130 50.030 ;
        RECT 122.970 50.030 123.260 76.860 ;
        RECT 123.750 59.270 124.150 79.010 ;
        RECT 123.450 58.770 124.150 59.270 ;
        RECT 124.550 50.030 124.840 76.850 ;
        RECT 122.970 49.030 124.840 50.030 ;
        RECT 126.680 50.030 126.970 76.860 ;
        RECT 127.450 59.270 127.850 79.010 ;
        RECT 127.170 58.770 127.850 59.270 ;
        RECT 128.260 50.030 128.550 76.850 ;
        RECT 126.680 49.030 128.550 50.030 ;
        RECT 130.390 50.030 130.680 76.860 ;
        RECT 131.150 59.270 131.550 79.010 ;
        RECT 130.900 58.770 131.550 59.270 ;
        RECT 131.970 50.030 132.260 76.850 ;
        RECT 130.390 49.030 132.260 50.030 ;
        RECT 134.100 50.030 134.390 76.860 ;
        RECT 134.850 59.270 135.250 79.010 ;
        RECT 134.570 58.770 135.250 59.270 ;
        RECT 135.680 50.030 135.970 76.850 ;
        RECT 134.100 49.030 135.970 50.030 ;
        RECT 80.925 39.985 81.430 40.375 ;
        RECT 74.370 38.690 74.880 39.080 ;
        RECT 71.375 35.150 71.880 37.790 ;
        RECT 74.375 37.400 74.875 38.690 ;
        RECT 80.925 37.790 81.425 39.985 ;
        RECT 83.925 39.080 84.425 42.950 ;
        RECT 98.600 42.350 99.500 42.800 ;
        RECT 99.900 42.350 100.800 42.800 ;
        RECT 101.200 42.350 102.100 42.800 ;
        RECT 102.500 42.350 103.400 42.800 ;
        RECT 90.475 39.980 90.980 40.370 ;
        RECT 90.475 39.080 90.975 39.980 ;
        RECT 83.920 38.690 84.430 39.080 ;
        RECT 90.475 38.690 90.980 39.080 ;
        RECT 80.925 35.150 81.430 37.790 ;
        RECT 83.925 37.400 84.425 38.690 ;
        RECT 90.475 37.790 90.975 38.690 ;
        RECT 90.475 35.150 90.980 37.790 ;
        RECT 92.250 37.450 92.750 41.950 ;
        RECT 103.550 35.150 104.050 48.700 ;
        RECT 108.590 48.040 109.600 49.020 ;
        RECT 112.280 48.050 113.290 49.030 ;
        RECT 116.010 48.060 117.000 49.030 ;
        RECT 108.590 46.940 111.400 48.040 ;
        RECT 112.280 46.950 114.890 48.050 ;
        RECT 116.010 46.960 118.410 48.060 ;
        RECT 119.700 48.050 120.720 49.030 ;
        RECT 123.410 48.070 124.410 49.030 ;
        RECT 127.130 48.080 128.140 49.030 ;
        RECT 112.280 46.940 114.880 46.950 ;
        RECT 119.700 46.940 121.920 48.050 ;
        RECT 123.410 46.960 125.430 48.070 ;
        RECT 127.130 46.950 128.910 48.080 ;
        RECT 130.840 48.060 131.840 49.030 ;
        RECT 130.840 46.950 132.420 48.060 ;
        RECT 132.810 46.460 134.560 48.060 ;
        RECT 134.940 46.960 135.940 49.030 ;
        RECT 132.810 45.300 137.720 46.460 ;
        RECT 132.810 44.800 134.560 45.300 ;
        RECT 20.050 19.100 20.550 21.200 ;
        RECT 21.050 19.600 21.550 30.350 ;
        RECT 21.900 23.680 22.400 32.400 ;
        RECT 26.040 23.680 26.540 32.350 ;
        RECT 29.040 21.600 29.540 30.600 ;
        RECT 35.680 23.680 36.180 32.400 ;
        RECT 38.680 20.600 39.180 30.600 ;
        RECT 45.320 23.680 45.820 32.400 ;
        RECT 20.050 18.600 21.600 19.100 ;
        RECT 21.100 5.600 21.600 18.600 ;
        RECT 21.900 5.600 22.400 20.500 ;
        RECT 27.700 5.600 28.200 18.200 ;
        RECT 32.700 5.600 33.200 20.200 ;
        RECT 48.320 19.600 48.820 30.600 ;
        RECT 54.960 23.680 55.460 32.400 ;
        RECT 49.350 19.150 49.850 20.200 ;
        RECT 57.960 19.600 58.460 30.600 ;
        RECT 64.600 23.680 65.100 32.400 ;
        RECT 67.600 20.600 68.100 30.600 ;
        RECT 74.240 23.680 74.740 32.400 ;
        RECT 77.240 21.600 77.740 30.600 ;
        RECT 81.350 23.675 81.850 32.400 ;
        RECT 82.200 22.150 82.700 30.300 ;
        RECT 83.650 29.100 84.150 32.400 ;
        RECT 80.700 21.650 82.700 22.150 ;
        RECT 48.250 18.650 49.850 19.150 ;
        RECT 43.250 5.600 43.750 18.200 ;
        RECT 48.250 5.600 48.750 18.650 ;
        RECT 58.800 5.600 59.300 18.200 ;
        RECT 63.800 5.600 64.300 20.200 ;
        RECT 74.350 5.600 74.850 20.500 ;
        RECT 79.350 5.600 79.850 21.200 ;
        RECT 80.700 19.600 81.200 21.650 ;
        RECT 84.950 20.600 85.450 30.700 ;
        RECT 86.150 21.400 86.650 26.100 ;
        RECT 93.950 23.150 94.450 30.200 ;
        RECT 97.200 26.900 97.500 27.500 ;
        RECT 97.650 24.550 98.150 25.150 ;
        RECT 98.450 21.400 98.950 30.200 ;
        RECT 99.350 21.600 99.850 30.250 ;
        RECT 100.250 21.400 100.750 30.570 ;
        RECT 102.240 21.400 102.740 30.570 ;
        RECT 89.900 5.600 90.400 18.200 ;
        RECT 94.900 5.600 95.400 20.200 ;
        RECT 103.240 18.600 103.740 30.550 ;
        RECT 105.790 21.400 106.290 30.570 ;
        RECT 106.790 21.600 107.290 30.550 ;
        RECT 109.340 21.400 109.840 30.570 ;
        RECT 110.340 21.600 110.840 30.550 ;
        RECT 112.890 21.400 113.390 30.570 ;
        RECT 113.890 27.280 114.390 30.550 ;
        RECT 113.885 26.890 114.390 27.280 ;
        RECT 105.450 5.600 105.950 18.200 ;
        RECT 110.450 5.600 110.950 20.200 ;
        RECT 113.890 18.600 114.390 26.890 ;
        RECT 116.000 21.400 116.500 30.570 ;
        RECT 116.800 21.600 117.300 30.250 ;
        RECT 118.450 21.400 118.950 30.400 ;
        RECT 121.000 5.600 121.500 18.200 ;
        RECT 126.000 5.600 126.500 20.200 ;
        RECT 130.800 17.600 131.300 30.400 ;
        RECT 132.300 5.600 132.800 20.500 ;
        RECT 133.100 5.600 133.600 21.200 ;
      LAYER met3 ;
        RECT 43.655 155.995 45.235 156.325 ;
        RECT 62.165 155.995 63.745 156.325 ;
        RECT 80.675 155.995 82.255 156.325 ;
        RECT 99.185 155.995 100.765 156.325 ;
        RECT 52.910 153.275 54.490 153.605 ;
        RECT 71.420 153.275 73.000 153.605 ;
        RECT 89.930 153.275 91.510 153.605 ;
        RECT 108.440 153.275 110.020 153.605 ;
        RECT 43.655 150.555 45.235 150.885 ;
        RECT 62.165 150.555 63.745 150.885 ;
        RECT 80.675 150.555 82.255 150.885 ;
        RECT 99.185 150.555 100.765 150.885 ;
        RECT 52.910 147.835 54.490 148.165 ;
        RECT 71.420 147.835 73.000 148.165 ;
        RECT 89.930 147.835 91.510 148.165 ;
        RECT 108.440 147.835 110.020 148.165 ;
        RECT 43.655 145.115 45.235 145.445 ;
        RECT 62.165 145.115 63.745 145.445 ;
        RECT 80.675 145.115 82.255 145.445 ;
        RECT 99.185 145.115 100.765 145.445 ;
        RECT 52.910 142.395 54.490 142.725 ;
        RECT 71.420 142.395 73.000 142.725 ;
        RECT 89.930 142.395 91.510 142.725 ;
        RECT 108.440 142.395 110.020 142.725 ;
        RECT 64.695 142.370 65.025 142.385 ;
        RECT 64.020 142.070 65.025 142.370 ;
        RECT 45.835 141.690 46.165 141.705 ;
        RECT 64.020 141.690 64.320 142.070 ;
        RECT 64.695 142.055 65.025 142.070 ;
        RECT 45.835 141.390 64.320 141.690 ;
        RECT 45.835 141.375 46.165 141.390 ;
        RECT 43.655 139.675 45.235 140.005 ;
        RECT 62.165 139.675 63.745 140.005 ;
        RECT 80.675 139.675 82.255 140.005 ;
        RECT 99.185 139.675 100.765 140.005 ;
        RECT 52.910 136.955 54.490 137.285 ;
        RECT 71.420 136.955 73.000 137.285 ;
        RECT 89.930 136.955 91.510 137.285 ;
        RECT 108.440 136.955 110.020 137.285 ;
        RECT 43.655 134.235 45.235 134.565 ;
        RECT 62.165 134.235 63.745 134.565 ;
        RECT 80.675 134.235 82.255 134.565 ;
        RECT 99.185 134.235 100.765 134.565 ;
        RECT 52.910 131.515 54.490 131.845 ;
        RECT 71.420 131.515 73.000 131.845 ;
        RECT 89.930 131.515 91.510 131.845 ;
        RECT 108.440 131.515 110.020 131.845 ;
        RECT 43.655 128.795 45.235 129.125 ;
        RECT 62.165 128.795 63.745 129.125 ;
        RECT 80.675 128.795 82.255 129.125 ;
        RECT 99.185 128.795 100.765 129.125 ;
        RECT 52.910 126.075 54.490 126.405 ;
        RECT 71.420 126.075 73.000 126.405 ;
        RECT 89.930 126.075 91.510 126.405 ;
        RECT 108.440 126.075 110.020 126.405 ;
        RECT 43.655 123.355 45.235 123.685 ;
        RECT 62.165 123.355 63.745 123.685 ;
        RECT 80.675 123.355 82.255 123.685 ;
        RECT 99.185 123.355 100.765 123.685 ;
        RECT 52.910 120.635 54.490 120.965 ;
        RECT 71.420 120.635 73.000 120.965 ;
        RECT 89.930 120.635 91.510 120.965 ;
        RECT 108.440 120.635 110.020 120.965 ;
        RECT 43.655 117.915 45.235 118.245 ;
        RECT 62.165 117.915 63.745 118.245 ;
        RECT 80.675 117.915 82.255 118.245 ;
        RECT 99.185 117.915 100.765 118.245 ;
        RECT 52.910 115.195 54.490 115.525 ;
        RECT 71.420 115.195 73.000 115.525 ;
        RECT 89.930 115.195 91.510 115.525 ;
        RECT 108.440 115.195 110.020 115.525 ;
        RECT 43.655 112.475 45.235 112.805 ;
        RECT 62.165 112.475 63.745 112.805 ;
        RECT 80.675 112.475 82.255 112.805 ;
        RECT 99.185 112.475 100.765 112.805 ;
        RECT 52.910 109.755 54.490 110.085 ;
        RECT 71.420 109.755 73.000 110.085 ;
        RECT 89.930 109.755 91.510 110.085 ;
        RECT 108.440 109.755 110.020 110.085 ;
        RECT 43.655 107.035 45.235 107.365 ;
        RECT 62.165 107.035 63.745 107.365 ;
        RECT 80.675 107.035 82.255 107.365 ;
        RECT 99.185 107.035 100.765 107.365 ;
        RECT 52.910 104.315 54.490 104.645 ;
        RECT 71.420 104.315 73.000 104.645 ;
        RECT 89.930 104.315 91.510 104.645 ;
        RECT 108.440 104.315 110.020 104.645 ;
        RECT 43.655 101.595 45.235 101.925 ;
        RECT 62.165 101.595 63.745 101.925 ;
        RECT 80.675 101.595 82.255 101.925 ;
        RECT 99.185 101.595 100.765 101.925 ;
        RECT 52.910 98.875 54.490 99.205 ;
        RECT 71.420 98.875 73.000 99.205 ;
        RECT 89.930 98.875 91.510 99.205 ;
        RECT 108.440 98.875 110.020 99.205 ;
        RECT 43.655 96.155 45.235 96.485 ;
        RECT 62.165 96.155 63.745 96.485 ;
        RECT 80.675 96.155 82.255 96.485 ;
        RECT 99.185 96.155 100.765 96.485 ;
        RECT 52.910 93.435 54.490 93.765 ;
        RECT 71.420 93.435 73.000 93.765 ;
        RECT 89.930 93.435 91.510 93.765 ;
        RECT 108.440 93.435 110.020 93.765 ;
        RECT 43.655 90.715 45.235 91.045 ;
        RECT 62.165 90.715 63.745 91.045 ;
        RECT 80.675 90.715 82.255 91.045 ;
        RECT 99.185 90.715 100.765 91.045 ;
        RECT 52.910 87.995 54.490 88.325 ;
        RECT 71.420 87.995 73.000 88.325 ;
        RECT 89.930 87.995 91.510 88.325 ;
        RECT 108.440 87.995 110.020 88.325 ;
        RECT 43.655 85.275 45.235 85.605 ;
        RECT 62.165 85.275 63.745 85.605 ;
        RECT 80.675 85.275 82.255 85.605 ;
        RECT 99.185 85.275 100.765 85.605 ;
        RECT 52.910 82.555 54.490 82.885 ;
        RECT 71.420 82.555 73.000 82.885 ;
        RECT 89.930 82.555 91.510 82.885 ;
        RECT 108.440 82.555 110.020 82.885 ;
        RECT 22.800 75.110 23.300 75.150 ;
        RECT 22.775 74.720 23.325 75.110 ;
        RECT 22.800 72.770 23.300 74.720 ;
        RECT 23.800 74.150 24.300 76.550 ;
        RECT 24.850 75.610 25.350 77.050 ;
        RECT 24.825 75.010 25.375 75.610 ;
        RECT 24.850 74.150 25.350 75.010 ;
        RECT 23.775 73.550 24.325 74.150 ;
        RECT 24.825 73.550 25.375 74.150 ;
        RECT 22.775 72.380 23.325 72.770 ;
        RECT 21.800 72.085 22.300 72.250 ;
        RECT 21.775 71.485 22.325 72.085 ;
        RECT 21.800 70.550 22.300 71.485 ;
        RECT 22.800 71.190 23.300 72.380 ;
        RECT 22.705 70.800 23.300 71.190 ;
        RECT 21.775 69.950 22.325 70.550 ;
        RECT 20.325 68.800 21.375 69.900 ;
        RECT 21.800 68.900 22.300 69.950 ;
        RECT 22.800 69.900 23.300 70.800 ;
        RECT 22.775 69.300 23.325 69.900 ;
        RECT 23.800 69.850 24.300 73.550 ;
        RECT 24.850 69.850 25.350 73.550 ;
        RECT 25.850 69.900 26.350 76.550 ;
        RECT 28.800 75.900 29.300 77.050 ;
        RECT 28.775 75.510 29.325 75.900 ;
        RECT 28.800 72.770 29.300 75.510 ;
        RECT 29.800 75.110 30.800 75.950 ;
        RECT 29.775 74.720 30.825 75.110 ;
        RECT 28.775 72.380 29.325 72.770 ;
        RECT 28.800 71.190 29.300 72.380 ;
        RECT 29.800 71.980 30.800 74.720 ;
        RECT 29.775 71.585 30.825 71.980 ;
        RECT 28.775 70.800 29.325 71.190 ;
        RECT 28.800 70.000 29.300 70.800 ;
        RECT 29.800 70.400 30.800 71.585 ;
        RECT 42.350 71.450 43.400 71.550 ;
        RECT 47.680 71.450 48.280 71.475 ;
        RECT 69.170 71.450 69.770 71.475 ;
        RECT 88.410 71.450 89.010 71.475 ;
        RECT 40.000 70.950 89.010 71.450 ;
        RECT 47.680 70.925 48.280 70.950 ;
        RECT 69.170 70.925 69.770 70.950 ;
        RECT 88.410 70.925 89.010 70.950 ;
        RECT 29.775 70.010 30.825 70.400 ;
        RECT 25.825 69.300 26.375 69.900 ;
        RECT 22.800 69.100 23.300 69.300 ;
        RECT 20.350 67.900 21.350 68.800 ;
        RECT 21.775 68.300 22.325 68.900 ;
        RECT 29.800 68.300 30.800 70.010 ;
        RECT 20.000 37.500 38.860 67.900 ;
        RECT 100.400 64.350 101.000 64.375 ;
        RECT 100.400 63.850 104.800 64.350 ;
        RECT 100.400 63.825 101.000 63.850 ;
        RECT 62.280 59.950 62.885 59.975 ;
        RECT 76.060 59.950 76.660 59.975 ;
        RECT 97.700 59.950 98.300 59.975 ;
        RECT 99.490 59.950 99.880 59.975 ;
        RECT 102.070 59.950 102.460 59.975 ;
        RECT 48.400 59.450 103.750 59.950 ;
        RECT 62.280 59.425 62.885 59.450 ;
        RECT 76.060 59.425 76.660 59.450 ;
        RECT 97.700 59.425 98.300 59.450 ;
        RECT 99.490 59.425 99.880 59.450 ;
        RECT 102.070 59.425 102.460 59.450 ;
        RECT 47.550 58.950 48.150 58.975 ;
        RECT 55.390 58.950 55.990 58.975 ;
        RECT 82.950 58.950 83.550 58.975 ;
        RECT 88.550 58.950 89.150 58.975 ;
        RECT 40.700 58.450 95.700 58.950 ;
        RECT 47.550 58.425 48.150 58.450 ;
        RECT 55.390 58.425 55.990 58.450 ;
        RECT 82.950 58.425 83.550 58.450 ;
        RECT 88.550 58.425 89.150 58.450 ;
        RECT 68.550 57.950 69.150 57.975 ;
        RECT 40.000 57.450 95.700 57.950 ;
        RECT 68.550 57.425 69.150 57.450 ;
        RECT 67.550 56.950 68.150 56.975 ;
        RECT 40.000 56.450 95.700 56.950 ;
        RECT 67.550 56.425 68.150 56.450 ;
        RECT 98.200 49.250 98.590 49.275 ;
        RECT 100.780 49.250 101.170 49.275 ;
        RECT 103.360 49.250 103.750 49.275 ;
        RECT 98.200 48.750 103.900 49.250 ;
        RECT 98.200 48.725 98.590 48.750 ;
        RECT 100.780 48.725 101.170 48.750 ;
        RECT 103.360 48.725 103.750 48.750 ;
        RECT 55.225 42.900 55.825 42.925 ;
        RECT 60.050 42.900 60.650 42.925 ;
        RECT 82.300 42.900 82.900 42.925 ;
        RECT 83.875 42.900 84.475 42.925 ;
        RECT 41.100 42.400 103.700 42.900 ;
        RECT 55.225 42.375 55.825 42.400 ;
        RECT 60.050 42.375 60.650 42.400 ;
        RECT 82.300 42.375 82.900 42.400 ;
        RECT 83.875 42.375 84.475 42.400 ;
        RECT 98.550 42.375 99.550 42.400 ;
        RECT 99.850 42.375 100.850 42.400 ;
        RECT 101.150 42.375 102.150 42.400 ;
        RECT 102.450 42.375 103.450 42.400 ;
        RECT 43.900 41.900 44.500 41.925 ;
        RECT 53.800 41.900 54.400 41.925 ;
        RECT 64.775 41.900 65.375 41.925 ;
        RECT 74.325 41.900 74.925 41.925 ;
        RECT 76.050 41.900 76.650 41.925 ;
        RECT 92.200 41.900 92.800 41.925 ;
        RECT 41.100 41.400 95.600 41.900 ;
        RECT 43.900 41.375 44.500 41.400 ;
        RECT 53.800 41.375 54.400 41.400 ;
        RECT 64.775 41.375 65.375 41.400 ;
        RECT 74.325 41.375 74.925 41.400 ;
        RECT 76.050 41.375 76.650 41.400 ;
        RECT 92.200 41.375 92.800 41.400 ;
        RECT 29.800 35.000 30.800 37.100 ;
        RECT 97.150 27.450 97.550 27.475 ;
        RECT 82.300 27.425 97.550 27.450 ;
        RECT 82.150 26.950 97.550 27.425 ;
        RECT 82.150 26.875 82.750 26.950 ;
        RECT 97.150 26.925 97.550 26.950 ;
        RECT 93.900 25.100 94.500 25.125 ;
        RECT 97.600 25.100 98.200 25.125 ;
        RECT 93.900 24.600 98.650 25.100 ;
        RECT 93.900 24.575 94.500 24.600 ;
        RECT 97.600 24.575 98.200 24.600 ;
        RECT 28.990 22.150 29.590 22.175 ;
        RECT 77.190 22.150 77.790 22.175 ;
        RECT 99.300 22.150 99.900 22.175 ;
        RECT 106.740 22.150 107.340 22.175 ;
        RECT 110.290 22.150 110.890 22.175 ;
        RECT 116.750 22.150 117.350 22.175 ;
        RECT 21.750 21.650 132.950 22.150 ;
        RECT 28.990 21.625 29.590 21.650 ;
        RECT 77.190 21.625 77.790 21.650 ;
        RECT 99.300 21.625 99.900 21.650 ;
        RECT 106.740 21.625 107.340 21.650 ;
        RECT 110.290 21.625 110.890 21.650 ;
        RECT 116.750 21.625 117.350 21.650 ;
        RECT 20.000 21.150 20.600 21.175 ;
        RECT 38.630 21.150 39.230 21.175 ;
        RECT 67.550 21.150 68.150 21.175 ;
        RECT 79.300 21.150 79.900 21.175 ;
        RECT 84.900 21.150 85.500 21.175 ;
        RECT 133.050 21.150 133.650 21.175 ;
        RECT 20.000 20.650 133.650 21.150 ;
        RECT 20.000 20.625 20.600 20.650 ;
        RECT 38.630 20.625 39.230 20.650 ;
        RECT 67.550 20.625 68.150 20.650 ;
        RECT 79.300 20.625 79.900 20.650 ;
        RECT 84.900 20.625 85.500 20.650 ;
        RECT 133.050 20.625 133.650 20.650 ;
        RECT 21.000 20.150 21.600 20.175 ;
        RECT 32.650 20.150 33.250 20.175 ;
        RECT 48.270 20.150 48.870 20.175 ;
        RECT 49.300 20.150 49.900 20.175 ;
        RECT 57.910 20.150 58.510 20.175 ;
        RECT 63.750 20.150 64.350 20.175 ;
        RECT 80.650 20.150 81.250 20.175 ;
        RECT 94.850 20.150 95.450 20.175 ;
        RECT 110.400 20.150 111.000 20.175 ;
        RECT 125.950 20.150 126.550 20.175 ;
        RECT 21.000 19.650 132.950 20.150 ;
        RECT 21.000 19.625 21.600 19.650 ;
        RECT 32.650 19.625 33.250 19.650 ;
        RECT 48.270 19.625 48.870 19.650 ;
        RECT 49.300 19.625 49.900 19.650 ;
        RECT 57.910 19.625 58.510 19.650 ;
        RECT 63.750 19.625 64.350 19.650 ;
        RECT 80.650 19.625 81.250 19.650 ;
        RECT 94.850 19.625 95.450 19.650 ;
        RECT 110.400 19.625 111.000 19.650 ;
        RECT 125.950 19.625 126.550 19.650 ;
        RECT 103.190 19.150 103.790 19.175 ;
        RECT 113.840 19.150 114.440 19.175 ;
        RECT 21.750 18.650 134.250 19.150 ;
        RECT 103.190 18.625 103.790 18.650 ;
        RECT 113.840 18.625 114.440 18.650 ;
        RECT 27.650 18.150 28.250 18.175 ;
        RECT 43.200 18.150 43.800 18.175 ;
        RECT 58.750 18.150 59.350 18.175 ;
        RECT 89.850 18.150 90.450 18.175 ;
        RECT 105.400 18.150 106.000 18.175 ;
        RECT 120.950 18.150 121.550 18.175 ;
        RECT 130.750 18.150 131.350 18.175 ;
        RECT 21.750 17.650 132.950 18.150 ;
        RECT 27.650 17.625 28.250 17.650 ;
        RECT 43.200 17.625 43.800 17.650 ;
        RECT 58.750 17.625 59.350 17.650 ;
        RECT 89.850 17.625 90.450 17.650 ;
        RECT 105.400 17.625 106.000 17.650 ;
        RECT 120.950 17.625 121.550 17.650 ;
        RECT 130.750 17.625 131.350 17.650 ;
      LAYER met4 ;
        RECT 43.645 82.480 45.245 156.400 ;
        RECT 52.900 82.480 54.500 156.400 ;
        RECT 62.155 82.480 63.755 156.400 ;
        RECT 71.410 82.480 73.010 156.400 ;
        RECT 80.665 82.480 82.265 156.400 ;
        RECT 89.920 82.480 91.520 156.400 ;
        RECT 99.175 82.480 100.775 156.400 ;
        RECT 108.430 82.480 110.030 156.400 ;
        RECT 106.205 77.205 107.815 78.425 ;
        RECT 29.795 68.345 30.805 68.855 ;
        RECT 29.800 67.505 30.800 68.345 ;
        RECT 20.395 37.895 37.005 67.505 ;
        RECT 29.800 37.055 30.800 37.895 ;
        RECT 38.360 37.560 38.840 67.840 ;
        RECT 29.795 36.045 30.805 37.055 ;
  END
END tt_um_cas_sensor_project
END LIBRARY

