** sch_path: /home/ttuser/test/inverter.sch
.subckt inverter VDD A Y VSS
*.PININFO VDD:I A:I Y:O VSS:I
XM2 Y A VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 m=1
XM1 Y A VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
.ends
.end
