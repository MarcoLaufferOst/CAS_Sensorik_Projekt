magic
tech sky130A
magscale 1 2
timestamp 1736976312
<< viali >>
rect 8585 15113 8619 15147
rect 1041 14909 1075 14943
rect 8493 14909 8527 14943
rect 1225 14773 1259 14807
rect 5273 14569 5307 14603
rect 6193 14569 6227 14603
rect 6561 14569 6595 14603
rect 4905 14501 4939 14535
rect 10701 14501 10735 14535
rect 4629 14433 4663 14467
rect 5365 14433 5399 14467
rect 6009 14433 6043 14467
rect 6285 14433 6319 14467
rect 6469 14433 6503 14467
rect 8769 14433 8803 14467
rect 10793 14433 10827 14467
rect 10977 14433 11011 14467
rect 12817 14433 12851 14467
rect 6745 14365 6779 14399
rect 7021 14365 7055 14399
rect 9045 14365 9079 14399
rect 11253 14365 11287 14399
rect 12725 14365 12759 14399
rect 5917 14229 5951 14263
rect 8493 14229 8527 14263
rect 10517 14229 10551 14263
rect 12909 14229 12943 14263
rect 4892 14025 4926 14059
rect 6377 14025 6411 14059
rect 7849 14025 7883 14059
rect 10425 14025 10459 14059
rect 11805 14025 11839 14059
rect 7297 13957 7331 13991
rect 10793 13957 10827 13991
rect 4629 13889 4663 13923
rect 6469 13889 6503 13923
rect 7665 13889 7699 13923
rect 8953 13889 8987 13923
rect 10977 13889 11011 13923
rect 7113 13821 7147 13855
rect 7205 13821 7239 13855
rect 7481 13821 7515 13855
rect 7757 13821 7791 13855
rect 9137 13821 9171 13855
rect 10517 13821 10551 13855
rect 10701 13821 10735 13855
rect 11713 13821 11747 13855
rect 8401 13685 8435 13719
rect 9321 13685 9355 13719
rect 10977 13685 11011 13719
rect 5273 13481 5307 13515
rect 7205 13481 7239 13515
rect 7941 13481 7975 13515
rect 8861 13481 8895 13515
rect 11529 13481 11563 13515
rect 8125 13413 8159 13447
rect 10425 13413 10459 13447
rect 10609 13413 10643 13447
rect 11161 13413 11195 13447
rect 3893 13345 3927 13379
rect 4813 13345 4847 13379
rect 5549 13345 5583 13379
rect 5641 13345 5675 13379
rect 7113 13345 7147 13379
rect 7389 13345 7423 13379
rect 7665 13345 7699 13379
rect 7849 13345 7883 13379
rect 8493 13345 8527 13379
rect 8585 13345 8619 13379
rect 8769 13345 8803 13379
rect 9045 13345 9079 13379
rect 9229 13345 9263 13379
rect 9505 13345 9539 13379
rect 9689 13345 9723 13379
rect 10149 13345 10183 13379
rect 10517 13345 10551 13379
rect 10701 13345 10735 13379
rect 10977 13345 11011 13379
rect 11253 13345 11287 13379
rect 11345 13345 11379 13379
rect 3065 13277 3099 13311
rect 4997 13277 5031 13311
rect 5181 13277 5215 13311
rect 6009 13277 6043 13311
rect 7021 13277 7055 13311
rect 7573 13277 7607 13311
rect 9321 13277 9355 13311
rect 9781 13277 9815 13311
rect 10425 13277 10459 13311
rect 6745 13209 6779 13243
rect 7481 13209 7515 13243
rect 8677 13209 8711 13243
rect 9137 13209 9171 13243
rect 10057 13209 10091 13243
rect 3801 13141 3835 13175
rect 4905 13141 4939 13175
rect 4997 13141 5031 13175
rect 5457 13141 5491 13175
rect 6653 13141 6687 13175
rect 6929 13141 6963 13175
rect 8125 13141 8159 13175
rect 9689 13141 9723 13175
rect 10241 13141 10275 13175
rect 4813 12937 4847 12971
rect 10057 12937 10091 12971
rect 12817 12937 12851 12971
rect 6285 12733 6319 12767
rect 8493 12733 8527 12767
rect 8953 12733 8987 12767
rect 9965 12733 9999 12767
rect 12725 12733 12759 12767
rect 6469 12665 6503 12699
rect 8217 12665 8251 12699
rect 8677 12665 8711 12699
rect 5641 12393 5675 12427
rect 6745 12393 6779 12427
rect 8217 12393 8251 12427
rect 8769 12393 8803 12427
rect 9781 12393 9815 12427
rect 12725 12393 12759 12427
rect 6469 12325 6503 12359
rect 8401 12325 8435 12359
rect 10195 12325 10229 12359
rect 10425 12325 10459 12359
rect 10701 12325 10735 12359
rect 11253 12325 11287 12359
rect 2053 12257 2087 12291
rect 3893 12257 3927 12291
rect 6009 12257 6043 12291
rect 6101 12257 6135 12291
rect 6377 12257 6411 12291
rect 6745 12257 6779 12291
rect 6929 12257 6963 12291
rect 7757 12257 7791 12291
rect 8309 12257 8343 12291
rect 8493 12257 8527 12291
rect 8677 12257 8711 12291
rect 9229 12257 9263 12291
rect 9505 12257 9539 12291
rect 10333 12257 10367 12291
rect 10517 12257 10551 12291
rect 2329 12189 2363 12223
rect 4169 12189 4203 12223
rect 10057 12189 10091 12223
rect 10977 12189 11011 12223
rect 5825 12121 5859 12155
rect 3801 12053 3835 12087
rect 8033 12053 8067 12087
rect 9321 12053 9355 12087
rect 4721 11849 4755 11883
rect 7665 11849 7699 11883
rect 12357 11849 12391 11883
rect 12633 11849 12667 11883
rect 14565 11849 14599 11883
rect 5641 11781 5675 11815
rect 9413 11781 9447 11815
rect 12265 11781 12299 11815
rect 6193 11713 6227 11747
rect 6745 11713 6779 11747
rect 12449 11713 12483 11747
rect 4629 11645 4663 11679
rect 5549 11645 5583 11679
rect 5733 11645 5767 11679
rect 5825 11645 5859 11679
rect 6009 11645 6043 11679
rect 6285 11645 6319 11679
rect 6561 11645 6595 11679
rect 6653 11645 6687 11679
rect 7297 11645 7331 11679
rect 7695 11645 7729 11679
rect 7849 11645 7883 11679
rect 8677 11645 8711 11679
rect 8861 11645 8895 11679
rect 9045 11645 9079 11679
rect 9321 11645 9355 11679
rect 9597 11645 9631 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 12541 11645 12575 11679
rect 14473 11645 14507 11679
rect 11437 11577 11471 11611
rect 5365 11509 5399 11543
rect 6469 11509 6503 11543
rect 8769 11509 8803 11543
rect 10885 11509 10919 11543
rect 5641 11305 5675 11339
rect 12725 11305 12759 11339
rect 5917 11237 5951 11271
rect 8217 11237 8251 11271
rect 8401 11237 8435 11271
rect 9413 11237 9447 11271
rect 10103 11237 10137 11271
rect 10333 11237 10367 11271
rect 10609 11237 10643 11271
rect 11253 11237 11287 11271
rect 3893 11169 3927 11203
rect 6009 11169 6043 11203
rect 6745 11169 6779 11203
rect 8309 11169 8343 11203
rect 8585 11169 8619 11203
rect 9045 11169 9079 11203
rect 9137 11169 9171 11203
rect 9689 11169 9723 11203
rect 9965 11169 9999 11203
rect 10241 11169 10275 11203
rect 10425 11169 10459 11203
rect 4169 11101 4203 11135
rect 7573 11101 7607 11135
rect 9321 11101 9355 11135
rect 9597 11101 9631 11135
rect 10977 11101 11011 11135
rect 6837 11033 6871 11067
rect 8769 10965 8803 10999
rect 9229 10965 9263 10999
rect 9413 10965 9447 10999
rect 9873 10965 9907 10999
rect 10885 10761 10919 10795
rect 11529 10761 11563 10795
rect 5825 10625 5859 10659
rect 7619 10625 7653 10659
rect 8953 10625 8987 10659
rect 6193 10557 6227 10591
rect 8217 10557 8251 10591
rect 9137 10557 9171 10591
rect 9505 10557 9539 10591
rect 11437 10557 11471 10591
rect 8125 10421 8159 10455
rect 8401 10421 8435 10455
rect 6285 10217 6319 10251
rect 10241 10217 10275 10251
rect 8769 10081 8803 10115
rect 9137 10081 9171 10115
rect 10333 10081 10367 10115
rect 6929 10013 6963 10047
rect 7389 9877 7423 9911
rect 6285 9605 6319 9639
rect 6469 9469 6503 9503
rect 6653 9469 6687 9503
rect 6745 9469 6779 9503
rect 8585 969 8619 1003
rect 8493 697 8527 731
<< metal1 >>
rect 552 15258 15364 15280
rect 552 15206 2249 15258
rect 2301 15206 2313 15258
rect 2365 15206 2377 15258
rect 2429 15206 2441 15258
rect 2493 15206 2505 15258
rect 2557 15206 5951 15258
rect 6003 15206 6015 15258
rect 6067 15206 6079 15258
rect 6131 15206 6143 15258
rect 6195 15206 6207 15258
rect 6259 15206 9653 15258
rect 9705 15206 9717 15258
rect 9769 15206 9781 15258
rect 9833 15206 9845 15258
rect 9897 15206 9909 15258
rect 9961 15206 13355 15258
rect 13407 15206 13419 15258
rect 13471 15206 13483 15258
rect 13535 15206 13547 15258
rect 13599 15206 13611 15258
rect 13663 15206 15364 15258
rect 552 15184 15364 15206
rect 8573 15147 8631 15153
rect 8573 15113 8585 15147
rect 8619 15144 8631 15147
rect 8754 15144 8760 15156
rect 8619 15116 8760 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 1026 14900 1032 14952
rect 1084 14900 1090 14952
rect 8478 14900 8484 14952
rect 8536 14900 8542 14952
rect 1213 14807 1271 14813
rect 1213 14773 1225 14807
rect 1259 14804 1271 14807
rect 3878 14804 3884 14816
rect 1259 14776 3884 14804
rect 1259 14773 1271 14776
rect 1213 14767 1271 14773
rect 3878 14764 3884 14776
rect 3936 14804 3942 14816
rect 4614 14804 4620 14816
rect 3936 14776 4620 14804
rect 3936 14764 3942 14776
rect 4614 14764 4620 14776
rect 4672 14764 4678 14816
rect 552 14714 15520 14736
rect 552 14662 4100 14714
rect 4152 14662 4164 14714
rect 4216 14662 4228 14714
rect 4280 14662 4292 14714
rect 4344 14662 4356 14714
rect 4408 14662 7802 14714
rect 7854 14662 7866 14714
rect 7918 14662 7930 14714
rect 7982 14662 7994 14714
rect 8046 14662 8058 14714
rect 8110 14662 11504 14714
rect 11556 14662 11568 14714
rect 11620 14662 11632 14714
rect 11684 14662 11696 14714
rect 11748 14662 11760 14714
rect 11812 14662 15206 14714
rect 15258 14662 15270 14714
rect 15322 14662 15334 14714
rect 15386 14662 15398 14714
rect 15450 14662 15462 14714
rect 15514 14662 15520 14714
rect 552 14640 15520 14662
rect 4430 14560 4436 14612
rect 4488 14600 4494 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 4488 14572 5273 14600
rect 4488 14560 4494 14572
rect 5261 14569 5273 14572
rect 5307 14569 5319 14603
rect 5261 14563 5319 14569
rect 5626 14560 5632 14612
rect 5684 14600 5690 14612
rect 6181 14603 6239 14609
rect 6181 14600 6193 14603
rect 5684 14572 6193 14600
rect 5684 14560 5690 14572
rect 6181 14569 6193 14572
rect 6227 14569 6239 14603
rect 6181 14563 6239 14569
rect 6549 14603 6607 14609
rect 6549 14569 6561 14603
rect 6595 14600 6607 14603
rect 7190 14600 7196 14612
rect 6595 14572 7196 14600
rect 6595 14569 6607 14572
rect 6549 14563 6607 14569
rect 7190 14560 7196 14572
rect 7248 14560 7254 14612
rect 8772 14572 11008 14600
rect 4893 14535 4951 14541
rect 4893 14501 4905 14535
rect 4939 14532 4951 14535
rect 7098 14532 7104 14544
rect 4939 14504 7104 14532
rect 4939 14501 4951 14504
rect 4893 14495 4951 14501
rect 4614 14424 4620 14476
rect 4672 14424 4678 14476
rect 5353 14467 5411 14473
rect 5353 14433 5365 14467
rect 5399 14464 5411 14467
rect 5810 14464 5816 14476
rect 5399 14436 5816 14464
rect 5399 14433 5411 14436
rect 5353 14427 5411 14433
rect 5810 14424 5816 14436
rect 5868 14424 5874 14476
rect 6012 14473 6040 14504
rect 7098 14492 7104 14504
rect 7156 14492 7162 14544
rect 7742 14492 7748 14544
rect 7800 14492 7806 14544
rect 5997 14467 6055 14473
rect 5997 14433 6009 14467
rect 6043 14433 6055 14467
rect 5997 14427 6055 14433
rect 6270 14424 6276 14476
rect 6328 14424 6334 14476
rect 6362 14424 6368 14476
rect 6420 14464 6426 14476
rect 8772 14473 8800 14572
rect 10689 14535 10747 14541
rect 10689 14532 10701 14535
rect 10258 14504 10701 14532
rect 10689 14501 10701 14504
rect 10735 14501 10747 14535
rect 10689 14495 10747 14501
rect 10980 14476 11008 14572
rect 11790 14492 11796 14544
rect 11848 14492 11854 14544
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 6420 14436 6469 14464
rect 6420 14424 6426 14436
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 8757 14467 8815 14473
rect 8757 14433 8769 14467
rect 8803 14433 8815 14467
rect 10778 14464 10784 14476
rect 8757 14427 8815 14433
rect 10244 14436 10784 14464
rect 4890 14356 4896 14408
rect 4948 14396 4954 14408
rect 6733 14399 6791 14405
rect 6733 14396 6745 14399
rect 4948 14368 6745 14396
rect 4948 14356 4954 14368
rect 6733 14365 6745 14368
rect 6779 14365 6791 14399
rect 6733 14359 6791 14365
rect 7006 14356 7012 14408
rect 7064 14356 7070 14408
rect 9030 14356 9036 14408
rect 9088 14356 9094 14408
rect 8202 14288 8208 14340
rect 8260 14328 8266 14340
rect 8260 14300 8892 14328
rect 8260 14288 8266 14300
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 5905 14263 5963 14269
rect 5905 14260 5917 14263
rect 5684 14232 5917 14260
rect 5684 14220 5690 14232
rect 5905 14229 5917 14232
rect 5951 14229 5963 14263
rect 5905 14223 5963 14229
rect 8478 14220 8484 14272
rect 8536 14220 8542 14272
rect 8864 14260 8892 14300
rect 10244 14260 10272 14436
rect 10778 14424 10784 14436
rect 10836 14424 10842 14476
rect 10962 14424 10968 14476
rect 11020 14424 11026 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12728 14436 12817 14464
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 12728 14405 12756 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14365 12771 14399
rect 12713 14359 12771 14365
rect 8864 14232 10272 14260
rect 10502 14220 10508 14272
rect 10560 14220 10566 14272
rect 12342 14220 12348 14272
rect 12400 14260 12406 14272
rect 12897 14263 12955 14269
rect 12897 14260 12909 14263
rect 12400 14232 12909 14260
rect 12400 14220 12406 14232
rect 12897 14229 12909 14232
rect 12943 14229 12955 14263
rect 12897 14223 12955 14229
rect 552 14170 15364 14192
rect 552 14118 2249 14170
rect 2301 14118 2313 14170
rect 2365 14118 2377 14170
rect 2429 14118 2441 14170
rect 2493 14118 2505 14170
rect 2557 14118 5951 14170
rect 6003 14118 6015 14170
rect 6067 14118 6079 14170
rect 6131 14118 6143 14170
rect 6195 14118 6207 14170
rect 6259 14118 9653 14170
rect 9705 14118 9717 14170
rect 9769 14118 9781 14170
rect 9833 14118 9845 14170
rect 9897 14118 9909 14170
rect 9961 14118 13355 14170
rect 13407 14118 13419 14170
rect 13471 14118 13483 14170
rect 13535 14118 13547 14170
rect 13599 14118 13611 14170
rect 13663 14118 15364 14170
rect 552 14096 15364 14118
rect 4880 14059 4938 14065
rect 4880 14025 4892 14059
rect 4926 14056 4938 14059
rect 4926 14028 5948 14056
rect 4926 14025 4938 14028
rect 4880 14019 4938 14025
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 4890 13920 4896 13932
rect 4663 13892 4896 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 5920 13920 5948 14028
rect 6362 14016 6368 14068
rect 6420 14016 6426 14068
rect 7098 14016 7104 14068
rect 7156 14056 7162 14068
rect 7156 14028 7696 14056
rect 7156 14016 7162 14028
rect 6380 13920 6408 14016
rect 6546 13948 6552 14000
rect 6604 13988 6610 14000
rect 7285 13991 7343 13997
rect 7285 13988 7297 13991
rect 6604 13960 7297 13988
rect 6604 13948 6610 13960
rect 7285 13957 7297 13960
rect 7331 13957 7343 13991
rect 7668 13988 7696 14028
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 7837 14059 7895 14065
rect 7837 14056 7849 14059
rect 7800 14028 7849 14056
rect 7800 14016 7806 14028
rect 7837 14025 7849 14028
rect 7883 14025 7895 14059
rect 7837 14019 7895 14025
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 10413 14059 10471 14065
rect 10413 14056 10425 14059
rect 10376 14028 10425 14056
rect 10376 14016 10382 14028
rect 10413 14025 10425 14028
rect 10459 14025 10471 14059
rect 10413 14019 10471 14025
rect 11790 14016 11796 14068
rect 11848 14016 11854 14068
rect 8202 13988 8208 14000
rect 7668 13960 8208 13988
rect 7285 13951 7343 13957
rect 6457 13923 6515 13929
rect 6457 13920 6469 13923
rect 5920 13892 6316 13920
rect 6380 13892 6469 13920
rect 6288 13852 6316 13892
rect 6457 13889 6469 13892
rect 6503 13889 6515 13923
rect 7653 13923 7711 13929
rect 7653 13920 7665 13923
rect 6457 13883 6515 13889
rect 6886 13892 7665 13920
rect 6886 13852 6914 13892
rect 7653 13889 7665 13892
rect 7699 13889 7711 13923
rect 7653 13883 7711 13889
rect 7760 13861 7788 13960
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 10686 13948 10692 14000
rect 10744 13988 10750 14000
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 10744 13960 10793 13988
rect 10744 13948 10750 13960
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 8478 13880 8484 13932
rect 8536 13920 8542 13932
rect 8941 13923 8999 13929
rect 8941 13920 8953 13923
rect 8536 13892 8953 13920
rect 8536 13880 8542 13892
rect 8941 13889 8953 13892
rect 8987 13889 8999 13923
rect 8941 13883 8999 13889
rect 10965 13923 11023 13929
rect 10965 13889 10977 13923
rect 11011 13920 11023 13923
rect 12342 13920 12348 13932
rect 11011 13892 12348 13920
rect 11011 13889 11023 13892
rect 10965 13883 11023 13889
rect 12342 13880 12348 13892
rect 12400 13880 12406 13932
rect 6288 13824 6914 13852
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7193 13855 7251 13861
rect 7193 13852 7205 13855
rect 7147 13824 7205 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7193 13821 7205 13824
rect 7239 13821 7251 13855
rect 7469 13855 7527 13861
rect 7469 13852 7481 13855
rect 7193 13815 7251 13821
rect 7300 13824 7481 13852
rect 5626 13744 5632 13796
rect 5684 13744 5690 13796
rect 6178 13744 6184 13796
rect 6236 13784 6242 13796
rect 7300 13784 7328 13824
rect 7469 13821 7481 13824
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 7745 13855 7803 13861
rect 7745 13821 7757 13855
rect 7791 13821 7803 13855
rect 7745 13815 7803 13821
rect 8202 13812 8208 13864
rect 8260 13852 8266 13864
rect 9125 13855 9183 13861
rect 9125 13852 9137 13855
rect 8260 13824 9137 13852
rect 8260 13812 8266 13824
rect 9125 13821 9137 13824
rect 9171 13821 9183 13855
rect 9125 13815 9183 13821
rect 10502 13812 10508 13864
rect 10560 13812 10566 13864
rect 10689 13855 10747 13861
rect 10689 13821 10701 13855
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 9214 13784 9220 13796
rect 6236 13756 7328 13784
rect 7392 13756 9220 13784
rect 6236 13744 6242 13756
rect 5534 13676 5540 13728
rect 5592 13716 5598 13728
rect 6914 13716 6920 13728
rect 5592 13688 6920 13716
rect 5592 13676 5598 13688
rect 6914 13676 6920 13688
rect 6972 13716 6978 13728
rect 7392 13716 7420 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9858 13744 9864 13796
rect 9916 13784 9922 13796
rect 10704 13784 10732 13815
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 10836 13824 11713 13852
rect 10836 13812 10842 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11701 13815 11759 13821
rect 9916 13756 10732 13784
rect 9916 13744 9922 13756
rect 6972 13688 7420 13716
rect 6972 13676 6978 13688
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 8389 13719 8447 13725
rect 8389 13716 8401 13719
rect 7708 13688 8401 13716
rect 7708 13676 7714 13688
rect 8389 13685 8401 13688
rect 8435 13685 8447 13719
rect 8389 13679 8447 13685
rect 8478 13676 8484 13728
rect 8536 13716 8542 13728
rect 9309 13719 9367 13725
rect 9309 13716 9321 13719
rect 8536 13688 9321 13716
rect 8536 13676 8542 13688
rect 9309 13685 9321 13688
rect 9355 13685 9367 13719
rect 9309 13679 9367 13685
rect 10965 13719 11023 13725
rect 10965 13685 10977 13719
rect 11011 13716 11023 13719
rect 11330 13716 11336 13728
rect 11011 13688 11336 13716
rect 11011 13685 11023 13688
rect 10965 13679 11023 13685
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 552 13626 15520 13648
rect 552 13574 4100 13626
rect 4152 13574 4164 13626
rect 4216 13574 4228 13626
rect 4280 13574 4292 13626
rect 4344 13574 4356 13626
rect 4408 13574 7802 13626
rect 7854 13574 7866 13626
rect 7918 13574 7930 13626
rect 7982 13574 7994 13626
rect 8046 13574 8058 13626
rect 8110 13574 11504 13626
rect 11556 13574 11568 13626
rect 11620 13574 11632 13626
rect 11684 13574 11696 13626
rect 11748 13574 11760 13626
rect 11812 13574 15206 13626
rect 15258 13574 15270 13626
rect 15322 13574 15334 13626
rect 15386 13574 15398 13626
rect 15450 13574 15462 13626
rect 15514 13574 15520 13626
rect 552 13552 15520 13574
rect 5261 13515 5319 13521
rect 5261 13481 5273 13515
rect 5307 13512 5319 13515
rect 6178 13512 6184 13524
rect 5307 13484 6184 13512
rect 5307 13481 5319 13484
rect 5261 13475 5319 13481
rect 6178 13472 6184 13484
rect 6236 13472 6242 13524
rect 7006 13472 7012 13524
rect 7064 13512 7070 13524
rect 7193 13515 7251 13521
rect 7193 13512 7205 13515
rect 7064 13484 7205 13512
rect 7064 13472 7070 13484
rect 7193 13481 7205 13484
rect 7239 13481 7251 13515
rect 7929 13515 7987 13521
rect 7929 13512 7941 13515
rect 7193 13475 7251 13481
rect 7852 13484 7941 13512
rect 5166 13404 5172 13456
rect 5224 13444 5230 13456
rect 5224 13416 7788 13444
rect 5224 13404 5230 13416
rect 3878 13336 3884 13388
rect 3936 13336 3942 13388
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13376 4859 13379
rect 4847 13348 5396 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 3050 13268 3056 13320
rect 3108 13268 3114 13320
rect 4982 13268 4988 13320
rect 5040 13268 5046 13320
rect 5166 13268 5172 13320
rect 5224 13268 5230 13320
rect 5368 13308 5396 13348
rect 5534 13336 5540 13388
rect 5592 13336 5598 13388
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 5675 13348 6316 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 5718 13308 5724 13320
rect 5368 13280 5724 13308
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 5868 13280 6009 13308
rect 5868 13268 5874 13280
rect 5997 13277 6009 13280
rect 6043 13277 6055 13311
rect 6288 13308 6316 13348
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 7101 13379 7159 13385
rect 7101 13376 7113 13379
rect 6788 13348 7113 13376
rect 6788 13336 6794 13348
rect 7101 13345 7113 13348
rect 7147 13345 7159 13379
rect 7101 13339 7159 13345
rect 7190 13336 7196 13388
rect 7248 13376 7254 13388
rect 7377 13379 7435 13385
rect 7377 13376 7389 13379
rect 7248 13348 7389 13376
rect 7248 13336 7254 13348
rect 7377 13345 7389 13348
rect 7423 13345 7435 13379
rect 7377 13339 7435 13345
rect 7650 13336 7656 13388
rect 7708 13336 7714 13388
rect 6288 13280 6914 13308
rect 5997 13271 6055 13277
rect 6454 13240 6460 13252
rect 5000 13212 6460 13240
rect 3786 13132 3792 13184
rect 3844 13132 3850 13184
rect 4798 13132 4804 13184
rect 4856 13172 4862 13184
rect 5000 13181 5028 13212
rect 6454 13200 6460 13212
rect 6512 13200 6518 13252
rect 6546 13200 6552 13252
rect 6604 13240 6610 13252
rect 6733 13243 6791 13249
rect 6733 13240 6745 13243
rect 6604 13212 6745 13240
rect 6604 13200 6610 13212
rect 6733 13209 6745 13212
rect 6779 13209 6791 13243
rect 6886 13240 6914 13280
rect 7006 13268 7012 13320
rect 7064 13268 7070 13320
rect 7558 13268 7564 13320
rect 7616 13308 7622 13320
rect 7760 13308 7788 13416
rect 7852 13385 7880 13484
rect 7929 13481 7941 13484
rect 7975 13481 7987 13515
rect 7929 13475 7987 13481
rect 8849 13515 8907 13521
rect 8849 13481 8861 13515
rect 8895 13512 8907 13515
rect 9030 13512 9036 13524
rect 8895 13484 9036 13512
rect 8895 13481 8907 13484
rect 8849 13475 8907 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 10134 13512 10140 13524
rect 9140 13484 10140 13512
rect 8113 13447 8171 13453
rect 8113 13413 8125 13447
rect 8159 13444 8171 13447
rect 9140 13444 9168 13484
rect 10134 13472 10140 13484
rect 10192 13472 10198 13524
rect 11238 13472 11244 13524
rect 11296 13512 11302 13524
rect 11517 13515 11575 13521
rect 11517 13512 11529 13515
rect 11296 13484 11529 13512
rect 11296 13472 11302 13484
rect 11517 13481 11529 13484
rect 11563 13481 11575 13515
rect 11517 13475 11575 13481
rect 10413 13447 10471 13453
rect 10413 13444 10425 13447
rect 8159 13416 9168 13444
rect 9508 13416 10425 13444
rect 8159 13413 8171 13416
rect 8113 13407 8171 13413
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13345 7895 13379
rect 8481 13379 8539 13385
rect 8481 13376 8493 13379
rect 7837 13339 7895 13345
rect 8036 13348 8493 13376
rect 8036 13308 8064 13348
rect 8481 13345 8493 13348
rect 8527 13345 8539 13379
rect 8481 13339 8539 13345
rect 8570 13336 8576 13388
rect 8628 13336 8634 13388
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13345 8815 13379
rect 8757 13339 8815 13345
rect 9033 13379 9091 13385
rect 9033 13345 9045 13379
rect 9079 13376 9091 13379
rect 9122 13376 9128 13388
rect 9079 13348 9128 13376
rect 9079 13345 9091 13348
rect 9033 13339 9091 13345
rect 7616 13280 8064 13308
rect 7616 13268 7622 13280
rect 8386 13268 8392 13320
rect 8444 13308 8450 13320
rect 8772 13308 8800 13339
rect 9122 13336 9128 13348
rect 9180 13336 9186 13388
rect 9508 13385 9536 13416
rect 10413 13413 10425 13416
rect 10459 13413 10471 13447
rect 10413 13407 10471 13413
rect 10597 13447 10655 13453
rect 10597 13413 10609 13447
rect 10643 13444 10655 13447
rect 11149 13447 11207 13453
rect 11149 13444 11161 13447
rect 10643 13416 11161 13444
rect 10643 13413 10655 13416
rect 10597 13407 10655 13413
rect 11149 13413 11161 13416
rect 11195 13413 11207 13447
rect 11149 13407 11207 13413
rect 9217 13379 9275 13385
rect 9217 13345 9229 13379
rect 9263 13376 9275 13379
rect 9493 13379 9551 13385
rect 9263 13348 9444 13376
rect 9263 13345 9275 13348
rect 9217 13339 9275 13345
rect 8444 13280 8800 13308
rect 8444 13268 8450 13280
rect 9306 13268 9312 13320
rect 9364 13268 9370 13320
rect 9416 13308 9444 13348
rect 9493 13345 9505 13379
rect 9539 13345 9551 13379
rect 9493 13339 9551 13345
rect 9677 13379 9735 13385
rect 9677 13345 9689 13379
rect 9723 13376 9735 13379
rect 9950 13376 9956 13388
rect 9723 13348 9956 13376
rect 9723 13345 9735 13348
rect 9677 13339 9735 13345
rect 9692 13308 9720 13339
rect 9950 13336 9956 13348
rect 10008 13336 10014 13388
rect 10042 13336 10048 13388
rect 10100 13336 10106 13388
rect 10134 13336 10140 13388
rect 10192 13336 10198 13388
rect 10505 13379 10563 13385
rect 10505 13376 10517 13379
rect 10244 13348 10517 13376
rect 9416 13280 9720 13308
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 10060 13308 10088 13336
rect 10244 13308 10272 13348
rect 10505 13345 10517 13348
rect 10551 13345 10563 13379
rect 10505 13339 10563 13345
rect 10686 13336 10692 13388
rect 10744 13336 10750 13388
rect 10778 13336 10784 13388
rect 10836 13376 10842 13388
rect 10965 13379 11023 13385
rect 10965 13376 10977 13379
rect 10836 13348 10977 13376
rect 10836 13336 10842 13348
rect 10965 13345 10977 13348
rect 11011 13345 11023 13379
rect 10965 13339 11023 13345
rect 11241 13379 11299 13385
rect 11241 13345 11253 13379
rect 11287 13345 11299 13379
rect 11241 13339 11299 13345
rect 9815 13280 10272 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 10413 13311 10471 13317
rect 10413 13308 10425 13311
rect 10376 13280 10425 13308
rect 10376 13268 10382 13280
rect 10413 13277 10425 13280
rect 10459 13277 10471 13311
rect 10413 13271 10471 13277
rect 6886 13212 7052 13240
rect 6733 13203 6791 13209
rect 4893 13175 4951 13181
rect 4893 13172 4905 13175
rect 4856 13144 4905 13172
rect 4856 13132 4862 13144
rect 4893 13141 4905 13144
rect 4939 13141 4951 13175
rect 4893 13135 4951 13141
rect 4985 13175 5043 13181
rect 4985 13141 4997 13175
rect 5031 13141 5043 13175
rect 4985 13135 5043 13141
rect 5166 13132 5172 13184
rect 5224 13172 5230 13184
rect 5445 13175 5503 13181
rect 5445 13172 5457 13175
rect 5224 13144 5457 13172
rect 5224 13132 5230 13144
rect 5445 13141 5457 13144
rect 5491 13141 5503 13175
rect 5445 13135 5503 13141
rect 6638 13132 6644 13184
rect 6696 13132 6702 13184
rect 6914 13132 6920 13184
rect 6972 13132 6978 13184
rect 7024 13172 7052 13212
rect 7466 13200 7472 13252
rect 7524 13200 7530 13252
rect 8665 13243 8723 13249
rect 8665 13240 8677 13243
rect 7576 13212 8677 13240
rect 7576 13172 7604 13212
rect 8665 13209 8677 13212
rect 8711 13240 8723 13243
rect 9125 13243 9183 13249
rect 9125 13240 9137 13243
rect 8711 13212 9137 13240
rect 8711 13209 8723 13212
rect 8665 13203 8723 13209
rect 9125 13209 9137 13212
rect 9171 13240 9183 13243
rect 9858 13240 9864 13252
rect 9171 13212 9864 13240
rect 9171 13209 9183 13212
rect 9125 13203 9183 13209
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 10045 13243 10103 13249
rect 10045 13209 10057 13243
rect 10091 13240 10103 13243
rect 11256 13240 11284 13339
rect 11330 13336 11336 13388
rect 11388 13336 11394 13388
rect 10091 13212 11284 13240
rect 10091 13209 10103 13212
rect 10045 13203 10103 13209
rect 7024 13144 7604 13172
rect 7650 13132 7656 13184
rect 7708 13172 7714 13184
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 7708 13144 8125 13172
rect 7708 13132 7714 13144
rect 8113 13141 8125 13144
rect 8159 13172 8171 13175
rect 8202 13172 8208 13184
rect 8159 13144 8208 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 9677 13175 9735 13181
rect 9677 13172 9689 13175
rect 9272 13144 9689 13172
rect 9272 13132 9278 13144
rect 9677 13141 9689 13144
rect 9723 13141 9735 13175
rect 9677 13135 9735 13141
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 10226 13172 10232 13184
rect 10008 13144 10232 13172
rect 10008 13132 10014 13144
rect 10226 13132 10232 13144
rect 10284 13172 10290 13184
rect 10686 13172 10692 13184
rect 10284 13144 10692 13172
rect 10284 13132 10290 13144
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 552 13082 15364 13104
rect 552 13030 2249 13082
rect 2301 13030 2313 13082
rect 2365 13030 2377 13082
rect 2429 13030 2441 13082
rect 2493 13030 2505 13082
rect 2557 13030 5951 13082
rect 6003 13030 6015 13082
rect 6067 13030 6079 13082
rect 6131 13030 6143 13082
rect 6195 13030 6207 13082
rect 6259 13030 9653 13082
rect 9705 13030 9717 13082
rect 9769 13030 9781 13082
rect 9833 13030 9845 13082
rect 9897 13030 9909 13082
rect 9961 13030 13355 13082
rect 13407 13030 13419 13082
rect 13471 13030 13483 13082
rect 13535 13030 13547 13082
rect 13599 13030 13611 13082
rect 13663 13030 15364 13082
rect 552 13008 15364 13030
rect 4801 12971 4859 12977
rect 4801 12937 4813 12971
rect 4847 12968 4859 12971
rect 4890 12968 4896 12980
rect 4847 12940 4896 12968
rect 4847 12937 4859 12940
rect 4801 12931 4859 12937
rect 4890 12928 4896 12940
rect 4948 12928 4954 12980
rect 4982 12928 4988 12980
rect 5040 12968 5046 12980
rect 6086 12968 6092 12980
rect 5040 12940 6092 12968
rect 5040 12928 5046 12940
rect 6086 12928 6092 12940
rect 6144 12928 6150 12980
rect 7006 12928 7012 12980
rect 7064 12968 7070 12980
rect 8754 12968 8760 12980
rect 7064 12940 8760 12968
rect 7064 12928 7070 12940
rect 8754 12928 8760 12940
rect 8812 12928 8818 12980
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10410 12968 10416 12980
rect 10091 12940 10416 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10410 12928 10416 12940
rect 10468 12968 10474 12980
rect 10778 12968 10784 12980
rect 10468 12940 10784 12968
rect 10468 12928 10474 12940
rect 10778 12928 10784 12940
rect 10836 12928 10842 12980
rect 12805 12971 12863 12977
rect 12805 12937 12817 12971
rect 12851 12968 12863 12971
rect 13078 12968 13084 12980
rect 12851 12940 13084 12968
rect 12851 12937 12863 12940
rect 12805 12931 12863 12937
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 7466 12900 7472 12912
rect 6886 12872 7472 12900
rect 4798 12792 4804 12844
rect 4856 12832 4862 12844
rect 5626 12832 5632 12844
rect 4856 12804 5632 12832
rect 4856 12792 4862 12804
rect 5626 12792 5632 12804
rect 5684 12832 5690 12844
rect 6886 12832 6914 12872
rect 7466 12860 7472 12872
rect 7524 12900 7530 12912
rect 8478 12900 8484 12912
rect 7524 12872 8484 12900
rect 7524 12860 7530 12872
rect 8478 12860 8484 12872
rect 8536 12860 8542 12912
rect 5684 12804 6914 12832
rect 8496 12804 9996 12832
rect 5684 12792 5690 12804
rect 6273 12767 6331 12773
rect 6273 12733 6285 12767
rect 6319 12764 6331 12767
rect 6319 12736 6914 12764
rect 6319 12733 6331 12736
rect 6273 12727 6331 12733
rect 6454 12656 6460 12708
rect 6512 12656 6518 12708
rect 6886 12696 6914 12736
rect 8386 12724 8392 12776
rect 8444 12764 8450 12776
rect 8496 12773 8524 12804
rect 8481 12767 8539 12773
rect 8481 12764 8493 12767
rect 8444 12736 8493 12764
rect 8444 12724 8450 12736
rect 8481 12733 8493 12736
rect 8527 12733 8539 12767
rect 8481 12727 8539 12733
rect 8570 12724 8576 12776
rect 8628 12764 8634 12776
rect 8938 12764 8944 12776
rect 8628 12736 8944 12764
rect 8628 12724 8634 12736
rect 8938 12724 8944 12736
rect 8996 12764 9002 12776
rect 9674 12764 9680 12776
rect 8996 12736 9680 12764
rect 8996 12724 9002 12736
rect 9674 12724 9680 12736
rect 9732 12764 9738 12776
rect 9858 12764 9864 12776
rect 9732 12736 9864 12764
rect 9732 12724 9738 12736
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 9968 12773 9996 12804
rect 9953 12767 10011 12773
rect 9953 12733 9965 12767
rect 9999 12733 10011 12767
rect 9953 12727 10011 12733
rect 12710 12724 12716 12776
rect 12768 12724 12774 12776
rect 8202 12696 8208 12708
rect 6886 12668 8208 12696
rect 8202 12656 8208 12668
rect 8260 12656 8266 12708
rect 8665 12699 8723 12705
rect 8665 12665 8677 12699
rect 8711 12696 8723 12699
rect 10134 12696 10140 12708
rect 8711 12668 10140 12696
rect 8711 12665 8723 12668
rect 8665 12659 8723 12665
rect 6086 12588 6092 12640
rect 6144 12628 6150 12640
rect 8680 12628 8708 12659
rect 10134 12656 10140 12668
rect 10192 12656 10198 12708
rect 6144 12600 8708 12628
rect 6144 12588 6150 12600
rect 552 12538 15520 12560
rect 552 12486 4100 12538
rect 4152 12486 4164 12538
rect 4216 12486 4228 12538
rect 4280 12486 4292 12538
rect 4344 12486 4356 12538
rect 4408 12486 7802 12538
rect 7854 12486 7866 12538
rect 7918 12486 7930 12538
rect 7982 12486 7994 12538
rect 8046 12486 8058 12538
rect 8110 12486 11504 12538
rect 11556 12486 11568 12538
rect 11620 12486 11632 12538
rect 11684 12486 11696 12538
rect 11748 12486 11760 12538
rect 11812 12486 15206 12538
rect 15258 12486 15270 12538
rect 15322 12486 15334 12538
rect 15386 12486 15398 12538
rect 15450 12486 15462 12538
rect 15514 12486 15520 12538
rect 552 12464 15520 12486
rect 4890 12424 4896 12436
rect 2148 12396 3924 12424
rect 2148 12356 2176 12396
rect 3786 12356 3792 12368
rect 2056 12328 2176 12356
rect 3542 12328 3792 12356
rect 2056 12297 2084 12328
rect 3786 12316 3792 12328
rect 3844 12316 3850 12368
rect 3896 12356 3924 12396
rect 4448 12396 4896 12424
rect 4448 12368 4476 12396
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 5629 12427 5687 12433
rect 5629 12393 5641 12427
rect 5675 12424 5687 12427
rect 5810 12424 5816 12436
rect 5675 12396 5816 12424
rect 5675 12393 5687 12396
rect 5629 12387 5687 12393
rect 5810 12384 5816 12396
rect 5868 12384 5874 12436
rect 6730 12424 6736 12436
rect 6012 12396 6736 12424
rect 4430 12356 4436 12368
rect 3896 12328 4436 12356
rect 3896 12297 3924 12328
rect 4430 12316 4436 12328
rect 4488 12316 4494 12368
rect 4706 12316 4712 12368
rect 4764 12316 4770 12368
rect 5718 12316 5724 12368
rect 5776 12316 5782 12368
rect 2041 12291 2099 12297
rect 2041 12257 2053 12291
rect 2087 12257 2099 12291
rect 2041 12251 2099 12257
rect 3881 12291 3939 12297
rect 3881 12257 3893 12291
rect 3927 12257 3939 12291
rect 5736 12288 5764 12316
rect 5810 12288 5816 12300
rect 5736 12260 5816 12288
rect 3881 12251 3939 12257
rect 5810 12248 5816 12260
rect 5868 12288 5874 12300
rect 6012 12297 6040 12396
rect 6730 12384 6736 12396
rect 6788 12384 6794 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8205 12427 8263 12433
rect 8205 12424 8217 12427
rect 7708 12396 8217 12424
rect 7708 12384 7714 12396
rect 8205 12393 8217 12396
rect 8251 12393 8263 12427
rect 8478 12424 8484 12436
rect 8205 12387 8263 12393
rect 8312 12396 8484 12424
rect 6457 12359 6515 12365
rect 6457 12325 6469 12359
rect 6503 12356 6515 12359
rect 6546 12356 6552 12368
rect 6503 12328 6552 12356
rect 6503 12325 6515 12328
rect 6457 12319 6515 12325
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 5997 12291 6055 12297
rect 5997 12288 6009 12291
rect 5868 12260 6009 12288
rect 5868 12248 5874 12260
rect 5997 12257 6009 12260
rect 6043 12257 6055 12291
rect 5997 12251 6055 12257
rect 6086 12248 6092 12300
rect 6144 12248 6150 12300
rect 6365 12291 6423 12297
rect 6365 12257 6377 12291
rect 6411 12288 6423 12291
rect 6638 12288 6644 12300
rect 6411 12260 6644 12288
rect 6411 12257 6423 12260
rect 6365 12251 6423 12257
rect 6638 12248 6644 12260
rect 6696 12248 6702 12300
rect 6733 12291 6791 12297
rect 6733 12257 6745 12291
rect 6779 12257 6791 12291
rect 6733 12251 6791 12257
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12220 2375 12223
rect 3050 12220 3056 12232
rect 2363 12192 3056 12220
rect 2363 12189 2375 12192
rect 2317 12183 2375 12189
rect 3050 12180 3056 12192
rect 3108 12180 3114 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 6104 12220 6132 12248
rect 6546 12220 6552 12232
rect 4203 12192 5856 12220
rect 6104 12192 6552 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 5828 12161 5856 12192
rect 6546 12180 6552 12192
rect 6604 12180 6610 12232
rect 5813 12155 5871 12161
rect 5813 12121 5825 12155
rect 5859 12121 5871 12155
rect 5813 12115 5871 12121
rect 6362 12112 6368 12164
rect 6420 12152 6426 12164
rect 6748 12152 6776 12251
rect 6914 12248 6920 12300
rect 6972 12248 6978 12300
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7024 12260 7757 12288
rect 6420 12124 6776 12152
rect 6420 12112 6426 12124
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 7024 12084 7052 12260
rect 7745 12257 7757 12260
rect 7791 12288 7803 12291
rect 8202 12288 8208 12300
rect 7791 12260 8208 12288
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 8202 12248 8208 12260
rect 8260 12248 8266 12300
rect 8312 12297 8340 12396
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 8754 12384 8760 12436
rect 8812 12424 8818 12436
rect 9769 12427 9827 12433
rect 8812 12396 9536 12424
rect 8812 12384 8818 12396
rect 8389 12359 8447 12365
rect 8389 12325 8401 12359
rect 8435 12356 8447 12359
rect 8570 12356 8576 12368
rect 8435 12328 8576 12356
rect 8435 12325 8447 12328
rect 8389 12319 8447 12325
rect 8570 12316 8576 12328
rect 8628 12356 8634 12368
rect 9306 12356 9312 12368
rect 8628 12328 9312 12356
rect 8628 12316 8634 12328
rect 9306 12316 9312 12328
rect 9364 12316 9370 12368
rect 8297 12291 8355 12297
rect 8297 12257 8309 12291
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 8481 12291 8539 12297
rect 8481 12257 8493 12291
rect 8527 12257 8539 12291
rect 8481 12251 8539 12257
rect 8665 12291 8723 12297
rect 8665 12257 8677 12291
rect 8711 12288 8723 12291
rect 8938 12288 8944 12300
rect 8711 12260 8944 12288
rect 8711 12257 8723 12260
rect 8665 12251 8723 12257
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8496 12220 8524 12251
rect 7616 12192 8524 12220
rect 7616 12180 7622 12192
rect 8680 12152 8708 12251
rect 8938 12248 8944 12260
rect 8996 12248 9002 12300
rect 9508 12297 9536 12396
rect 9769 12393 9781 12427
rect 9815 12393 9827 12427
rect 9769 12387 9827 12393
rect 9784 12356 9812 12387
rect 12710 12384 12716 12436
rect 12768 12384 12774 12436
rect 10183 12359 10241 12365
rect 10183 12356 10195 12359
rect 9784 12328 10195 12356
rect 10183 12325 10195 12328
rect 10229 12325 10241 12359
rect 10183 12319 10241 12325
rect 10410 12316 10416 12368
rect 10468 12316 10474 12368
rect 10689 12359 10747 12365
rect 10689 12325 10701 12359
rect 10735 12356 10747 12359
rect 11241 12359 11299 12365
rect 11241 12356 11253 12359
rect 10735 12328 11253 12356
rect 10735 12325 10747 12328
rect 10689 12319 10747 12325
rect 11241 12325 11253 12328
rect 11287 12325 11299 12359
rect 11241 12319 11299 12325
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9493 12291 9551 12297
rect 9263 12260 9444 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 8128 12124 8708 12152
rect 9416 12152 9444 12260
rect 9493 12257 9505 12291
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10318 12288 10324 12300
rect 9732 12260 10324 12288
rect 9732 12248 9738 12260
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 10502 12248 10508 12300
rect 10560 12248 10566 12300
rect 12618 12288 12624 12300
rect 12374 12260 12624 12288
rect 12618 12248 12624 12260
rect 12676 12248 12682 12300
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 10962 12180 10968 12232
rect 11020 12180 11026 12232
rect 10502 12152 10508 12164
rect 9416 12124 10508 12152
rect 3835 12056 7052 12084
rect 8021 12087 8079 12093
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 8021 12053 8033 12087
rect 8067 12084 8079 12087
rect 8128 12084 8156 12124
rect 10502 12112 10508 12124
rect 10560 12112 10566 12164
rect 8067 12056 8156 12084
rect 8067 12053 8079 12056
rect 8021 12047 8079 12053
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8386 12084 8392 12096
rect 8260 12056 8392 12084
rect 8260 12044 8266 12056
rect 8386 12044 8392 12056
rect 8444 12044 8450 12096
rect 9306 12044 9312 12096
rect 9364 12044 9370 12096
rect 552 11994 15364 12016
rect 552 11942 2249 11994
rect 2301 11942 2313 11994
rect 2365 11942 2377 11994
rect 2429 11942 2441 11994
rect 2493 11942 2505 11994
rect 2557 11942 5951 11994
rect 6003 11942 6015 11994
rect 6067 11942 6079 11994
rect 6131 11942 6143 11994
rect 6195 11942 6207 11994
rect 6259 11942 9653 11994
rect 9705 11942 9717 11994
rect 9769 11942 9781 11994
rect 9833 11942 9845 11994
rect 9897 11942 9909 11994
rect 9961 11942 13355 11994
rect 13407 11942 13419 11994
rect 13471 11942 13483 11994
rect 13535 11942 13547 11994
rect 13599 11942 13611 11994
rect 13663 11942 15364 11994
rect 552 11920 15364 11942
rect 4706 11840 4712 11892
rect 4764 11840 4770 11892
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 7653 11883 7711 11889
rect 7653 11880 7665 11883
rect 7616 11852 7665 11880
rect 7616 11840 7622 11852
rect 7653 11849 7665 11852
rect 7699 11849 7711 11883
rect 7653 11843 7711 11849
rect 8294 11840 8300 11892
rect 8352 11880 8358 11892
rect 8352 11852 9168 11880
rect 8352 11840 8358 11852
rect 5629 11815 5687 11821
rect 5629 11781 5641 11815
rect 5675 11812 5687 11815
rect 5810 11812 5816 11824
rect 5675 11784 5816 11812
rect 5675 11781 5687 11784
rect 5629 11775 5687 11781
rect 5810 11772 5816 11784
rect 5868 11772 5874 11824
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6420 11784 7696 11812
rect 6420 11772 6426 11784
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6733 11747 6791 11753
rect 6733 11744 6745 11747
rect 6227 11716 6745 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 6733 11713 6745 11716
rect 6779 11713 6791 11747
rect 6733 11707 6791 11713
rect 7668 11744 7696 11784
rect 9140 11744 9168 11852
rect 10042 11840 10048 11892
rect 10100 11880 10106 11892
rect 12345 11883 12403 11889
rect 12345 11880 12357 11883
rect 10100 11852 12357 11880
rect 10100 11840 10106 11852
rect 12345 11849 12357 11852
rect 12391 11849 12403 11883
rect 12345 11843 12403 11849
rect 12618 11840 12624 11892
rect 12676 11840 12682 11892
rect 14553 11883 14611 11889
rect 14553 11849 14565 11883
rect 14599 11880 14611 11883
rect 15010 11880 15016 11892
rect 14599 11852 15016 11880
rect 14599 11849 14611 11852
rect 14553 11843 14611 11849
rect 15010 11840 15016 11852
rect 15068 11840 15074 11892
rect 9401 11815 9459 11821
rect 9401 11781 9413 11815
rect 9447 11812 9459 11815
rect 10226 11812 10232 11824
rect 9447 11784 10232 11812
rect 9447 11781 9459 11784
rect 9401 11775 9459 11781
rect 10226 11772 10232 11784
rect 10284 11812 10290 11824
rect 12253 11815 12311 11821
rect 12253 11812 12265 11815
rect 10284 11784 12265 11812
rect 10284 11772 10290 11784
rect 12253 11781 12265 11784
rect 12299 11781 12311 11815
rect 12253 11775 12311 11781
rect 12437 11747 12495 11753
rect 7668 11716 8984 11744
rect 9140 11716 9628 11744
rect 7668 11688 7696 11716
rect 4614 11636 4620 11688
rect 4672 11636 4678 11688
rect 5534 11636 5540 11688
rect 5592 11636 5598 11688
rect 5626 11636 5632 11688
rect 5684 11676 5690 11688
rect 5721 11679 5779 11685
rect 5721 11676 5733 11679
rect 5684 11648 5733 11676
rect 5684 11636 5690 11648
rect 5721 11645 5733 11648
rect 5767 11645 5779 11679
rect 5721 11639 5779 11645
rect 5813 11679 5871 11685
rect 5813 11645 5825 11679
rect 5859 11676 5871 11679
rect 5997 11679 6055 11685
rect 5997 11676 6009 11679
rect 5859 11648 6009 11676
rect 5859 11645 5871 11648
rect 5813 11639 5871 11645
rect 5997 11645 6009 11648
rect 6043 11645 6055 11679
rect 5997 11639 6055 11645
rect 6273 11679 6331 11685
rect 6273 11645 6285 11679
rect 6319 11676 6331 11679
rect 6362 11676 6368 11688
rect 6319 11648 6368 11676
rect 6319 11645 6331 11648
rect 6273 11639 6331 11645
rect 5736 11608 5764 11639
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 6546 11636 6552 11688
rect 6604 11636 6610 11688
rect 6638 11636 6644 11688
rect 6696 11636 6702 11688
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 6880 11648 7297 11676
rect 6880 11636 6886 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 7650 11636 7656 11688
rect 7708 11685 7714 11688
rect 8680 11685 8708 11716
rect 7708 11679 7741 11685
rect 7729 11645 7741 11679
rect 7708 11639 7741 11645
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11645 7895 11679
rect 7837 11639 7895 11645
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11645 8723 11679
rect 8665 11639 8723 11645
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11645 8907 11679
rect 8956 11678 8984 11716
rect 9600 11685 9628 11716
rect 12437 11713 12449 11747
rect 12483 11744 12495 11747
rect 13078 11744 13084 11756
rect 12483 11716 13084 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 13078 11704 13084 11716
rect 13136 11704 13142 11756
rect 9033 11679 9091 11685
rect 9033 11678 9045 11679
rect 8956 11650 9045 11678
rect 8849 11639 8907 11645
rect 9033 11645 9045 11650
rect 9079 11645 9091 11679
rect 9033 11639 9091 11645
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 7708 11636 7714 11639
rect 6656 11608 6684 11636
rect 7852 11608 7880 11639
rect 8864 11608 8892 11639
rect 9324 11608 9352 11639
rect 9398 11608 9404 11620
rect 5736 11580 6684 11608
rect 7392 11580 9404 11608
rect 7392 11552 7420 11580
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 9950 11568 9956 11620
rect 10008 11608 10014 11620
rect 11425 11611 11483 11617
rect 11425 11608 11437 11611
rect 10008 11580 11437 11608
rect 10008 11568 10014 11580
rect 11425 11577 11437 11580
rect 11471 11577 11483 11611
rect 12084 11608 12112 11639
rect 12158 11636 12164 11688
rect 12216 11636 12222 11688
rect 12526 11636 12532 11688
rect 12584 11636 12590 11688
rect 12710 11636 12716 11688
rect 12768 11676 12774 11688
rect 14461 11679 14519 11685
rect 14461 11676 14473 11679
rect 12768 11648 14473 11676
rect 12768 11636 12774 11648
rect 14461 11645 14473 11648
rect 14507 11645 14519 11679
rect 14461 11639 14519 11645
rect 12728 11608 12756 11636
rect 12084 11580 12756 11608
rect 11425 11571 11483 11577
rect 5350 11500 5356 11552
rect 5408 11500 5414 11552
rect 6457 11543 6515 11549
rect 6457 11509 6469 11543
rect 6503 11540 6515 11543
rect 6914 11540 6920 11552
rect 6503 11512 6920 11540
rect 6503 11509 6515 11512
rect 6457 11503 6515 11509
rect 6914 11500 6920 11512
rect 6972 11540 6978 11552
rect 7374 11540 7380 11552
rect 6972 11512 7380 11540
rect 6972 11500 6978 11512
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 8757 11543 8815 11549
rect 8757 11509 8769 11543
rect 8803 11540 8815 11543
rect 9122 11540 9128 11552
rect 8803 11512 9128 11540
rect 8803 11509 8815 11512
rect 8757 11503 8815 11509
rect 9122 11500 9128 11512
rect 9180 11540 9186 11552
rect 10502 11540 10508 11552
rect 9180 11512 10508 11540
rect 9180 11500 9186 11512
rect 10502 11500 10508 11512
rect 10560 11500 10566 11552
rect 10873 11543 10931 11549
rect 10873 11509 10885 11543
rect 10919 11540 10931 11543
rect 10962 11540 10968 11552
rect 10919 11512 10968 11540
rect 10919 11509 10931 11512
rect 10873 11503 10931 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 552 11450 15520 11472
rect 552 11398 4100 11450
rect 4152 11398 4164 11450
rect 4216 11398 4228 11450
rect 4280 11398 4292 11450
rect 4344 11398 4356 11450
rect 4408 11398 7802 11450
rect 7854 11398 7866 11450
rect 7918 11398 7930 11450
rect 7982 11398 7994 11450
rect 8046 11398 8058 11450
rect 8110 11398 11504 11450
rect 11556 11398 11568 11450
rect 11620 11398 11632 11450
rect 11684 11398 11696 11450
rect 11748 11398 11760 11450
rect 11812 11398 15206 11450
rect 15258 11398 15270 11450
rect 15322 11398 15334 11450
rect 15386 11398 15398 11450
rect 15450 11398 15462 11450
rect 15514 11398 15520 11450
rect 552 11376 15520 11398
rect 5629 11339 5687 11345
rect 5629 11305 5641 11339
rect 5675 11336 5687 11339
rect 6270 11336 6276 11348
rect 5675 11308 6276 11336
rect 5675 11305 5687 11308
rect 5629 11299 5687 11305
rect 6270 11296 6276 11308
rect 6328 11336 6334 11348
rect 6822 11336 6828 11348
rect 6328 11308 6828 11336
rect 6328 11296 6334 11308
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 12158 11336 12164 11348
rect 9088 11308 12164 11336
rect 9088 11296 9094 11308
rect 4154 11268 4160 11280
rect 3896 11240 4160 11268
rect 3896 11209 3924 11240
rect 4154 11228 4160 11240
rect 4212 11268 4218 11280
rect 4430 11268 4436 11280
rect 4212 11240 4436 11268
rect 4212 11228 4218 11240
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 5905 11271 5963 11277
rect 5905 11268 5917 11271
rect 5382 11240 5917 11268
rect 5905 11237 5917 11240
rect 5951 11237 5963 11271
rect 5905 11231 5963 11237
rect 8205 11271 8263 11277
rect 8205 11237 8217 11271
rect 8251 11268 8263 11271
rect 8389 11271 8447 11277
rect 8389 11268 8401 11271
rect 8251 11240 8401 11268
rect 8251 11237 8263 11240
rect 8205 11231 8263 11237
rect 8389 11237 8401 11240
rect 8435 11237 8447 11271
rect 8389 11231 8447 11237
rect 8662 11228 8668 11280
rect 8720 11268 8726 11280
rect 9306 11268 9312 11280
rect 8720 11240 9312 11268
rect 8720 11228 8726 11240
rect 9306 11228 9312 11240
rect 9364 11268 9370 11280
rect 9401 11271 9459 11277
rect 9401 11268 9413 11271
rect 9364 11240 9413 11268
rect 9364 11228 9370 11240
rect 9401 11237 9413 11240
rect 9447 11237 9459 11271
rect 9401 11231 9459 11237
rect 9858 11228 9864 11280
rect 9916 11268 9922 11280
rect 10336 11277 10364 11308
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 12710 11296 12716 11348
rect 12768 11296 12774 11348
rect 10091 11271 10149 11277
rect 10091 11268 10103 11271
rect 9916 11240 10103 11268
rect 9916 11228 9922 11240
rect 10091 11237 10103 11240
rect 10137 11237 10149 11271
rect 10091 11231 10149 11237
rect 10321 11271 10379 11277
rect 10321 11237 10333 11271
rect 10367 11237 10379 11271
rect 10321 11231 10379 11237
rect 10597 11271 10655 11277
rect 10597 11237 10609 11271
rect 10643 11268 10655 11271
rect 11241 11271 11299 11277
rect 11241 11268 11253 11271
rect 10643 11240 11253 11268
rect 10643 11237 10655 11240
rect 10597 11231 10655 11237
rect 11241 11237 11253 11240
rect 11287 11237 11299 11271
rect 11241 11231 11299 11237
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 11572 11240 11730 11268
rect 11572 11228 11578 11240
rect 3881 11203 3939 11209
rect 3881 11169 3893 11203
rect 3927 11169 3939 11203
rect 3881 11163 3939 11169
rect 5997 11203 6055 11209
rect 5997 11169 6009 11203
rect 6043 11200 6055 11203
rect 6733 11203 6791 11209
rect 6733 11200 6745 11203
rect 6043 11172 6745 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 6733 11169 6745 11172
rect 6779 11200 6791 11203
rect 7006 11200 7012 11212
rect 6779 11172 7012 11200
rect 6779 11169 6791 11172
rect 6733 11163 6791 11169
rect 7006 11160 7012 11172
rect 7064 11200 7070 11212
rect 7282 11200 7288 11212
rect 7064 11172 7288 11200
rect 7064 11160 7070 11172
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 5350 11132 5356 11144
rect 4203 11104 5356 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 5350 11092 5356 11104
rect 5408 11092 5414 11144
rect 7374 11092 7380 11144
rect 7432 11132 7438 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 7432 11104 7573 11132
rect 7432 11092 7438 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 8312 11132 8340 11163
rect 8570 11160 8576 11212
rect 8628 11160 8634 11212
rect 9030 11160 9036 11212
rect 9088 11160 9094 11212
rect 9122 11160 9128 11212
rect 9180 11160 9186 11212
rect 9490 11160 9496 11212
rect 9548 11198 9554 11212
rect 9677 11203 9735 11209
rect 9677 11200 9689 11203
rect 9600 11198 9689 11200
rect 9548 11172 9689 11198
rect 9548 11170 9628 11172
rect 9548 11160 9554 11170
rect 9677 11169 9689 11172
rect 9723 11169 9735 11203
rect 9677 11163 9735 11169
rect 9950 11160 9956 11212
rect 10008 11160 10014 11212
rect 10226 11160 10232 11212
rect 10284 11160 10290 11212
rect 10413 11203 10471 11209
rect 10413 11169 10425 11203
rect 10459 11200 10471 11203
rect 10502 11200 10508 11212
rect 10459 11172 10508 11200
rect 10459 11169 10471 11172
rect 10413 11163 10471 11169
rect 10502 11160 10508 11172
rect 10560 11160 10566 11212
rect 8478 11132 8484 11144
rect 8312 11104 8484 11132
rect 7561 11095 7619 11101
rect 8478 11092 8484 11104
rect 8536 11132 8542 11144
rect 9048 11132 9076 11160
rect 8536 11104 9076 11132
rect 9309 11135 9367 11141
rect 8536 11092 8542 11104
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9585 11135 9643 11141
rect 9585 11101 9597 11135
rect 9631 11132 9643 11135
rect 10042 11132 10048 11144
rect 9631 11104 10048 11132
rect 9631 11101 9643 11104
rect 9585 11095 9643 11101
rect 6825 11067 6883 11073
rect 6825 11033 6837 11067
rect 6871 11064 6883 11067
rect 6914 11064 6920 11076
rect 6871 11036 6920 11064
rect 6871 11033 6883 11036
rect 6825 11027 6883 11033
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 9324 11064 9352 11095
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10244 11064 10272 11160
rect 10962 11092 10968 11144
rect 11020 11092 11026 11144
rect 9324 11036 10272 11064
rect 8754 10956 8760 11008
rect 8812 10956 8818 11008
rect 9214 10956 9220 11008
rect 9272 10956 9278 11008
rect 9398 10956 9404 11008
rect 9456 10956 9462 11008
rect 9858 10956 9864 11008
rect 9916 10956 9922 11008
rect 552 10906 15364 10928
rect 552 10854 2249 10906
rect 2301 10854 2313 10906
rect 2365 10854 2377 10906
rect 2429 10854 2441 10906
rect 2493 10854 2505 10906
rect 2557 10854 5951 10906
rect 6003 10854 6015 10906
rect 6067 10854 6079 10906
rect 6131 10854 6143 10906
rect 6195 10854 6207 10906
rect 6259 10854 9653 10906
rect 9705 10854 9717 10906
rect 9769 10854 9781 10906
rect 9833 10854 9845 10906
rect 9897 10854 9909 10906
rect 9961 10854 13355 10906
rect 13407 10854 13419 10906
rect 13471 10854 13483 10906
rect 13535 10854 13547 10906
rect 13599 10854 13611 10906
rect 13663 10854 15364 10906
rect 552 10832 15364 10854
rect 9490 10792 9496 10804
rect 8956 10764 9496 10792
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 7650 10665 7656 10668
rect 5813 10659 5871 10665
rect 5813 10656 5825 10659
rect 4212 10628 5825 10656
rect 4212 10616 4218 10628
rect 5813 10625 5825 10628
rect 5859 10625 5871 10659
rect 7607 10659 7656 10665
rect 7607 10656 7619 10659
rect 7563 10628 7619 10656
rect 5813 10619 5871 10625
rect 7607 10625 7619 10628
rect 7653 10625 7656 10659
rect 7607 10619 7656 10625
rect 7650 10616 7656 10619
rect 7708 10656 7714 10668
rect 8956 10665 8984 10764
rect 9490 10752 9496 10764
rect 9548 10752 9554 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10318 10792 10324 10804
rect 10100 10764 10324 10792
rect 10100 10752 10106 10764
rect 10318 10752 10324 10764
rect 10376 10792 10382 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 10376 10764 10885 10792
rect 10376 10752 10382 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 11514 10752 11520 10804
rect 11572 10752 11578 10804
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 7708 10628 8953 10656
rect 7708 10616 7714 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 10962 10656 10968 10668
rect 8941 10619 8999 10625
rect 9140 10628 10968 10656
rect 9140 10600 9168 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6270 10588 6276 10600
rect 6227 10560 6276 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6270 10548 6276 10560
rect 6328 10548 6334 10600
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 8205 10591 8263 10597
rect 8205 10588 8217 10591
rect 7064 10560 8217 10588
rect 7064 10548 7070 10560
rect 8205 10557 8217 10560
rect 8251 10588 8263 10591
rect 8251 10560 8984 10588
rect 8251 10557 8263 10560
rect 8205 10551 8263 10557
rect 6914 10480 6920 10532
rect 6972 10480 6978 10532
rect 8113 10455 8171 10461
rect 8113 10421 8125 10455
rect 8159 10452 8171 10455
rect 8202 10452 8208 10464
rect 8159 10424 8208 10452
rect 8159 10421 8171 10424
rect 8113 10415 8171 10421
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8386 10412 8392 10464
rect 8444 10412 8450 10464
rect 8956 10452 8984 10560
rect 9122 10548 9128 10600
rect 9180 10548 9186 10600
rect 9214 10548 9220 10600
rect 9272 10588 9278 10600
rect 9493 10591 9551 10597
rect 9493 10588 9505 10591
rect 9272 10560 9505 10588
rect 9272 10548 9278 10560
rect 9493 10557 9505 10560
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 11425 10591 11483 10597
rect 11425 10588 11437 10591
rect 10376 10560 11437 10588
rect 10376 10548 10382 10560
rect 11425 10557 11437 10560
rect 11471 10588 11483 10591
rect 12526 10588 12532 10600
rect 11471 10560 12532 10588
rect 11471 10557 11483 10560
rect 11425 10551 11483 10557
rect 12526 10548 12532 10560
rect 12584 10548 12590 10600
rect 10226 10480 10232 10532
rect 10284 10480 10290 10532
rect 10318 10452 10324 10464
rect 8956 10424 10324 10452
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 552 10362 15520 10384
rect 552 10310 4100 10362
rect 4152 10310 4164 10362
rect 4216 10310 4228 10362
rect 4280 10310 4292 10362
rect 4344 10310 4356 10362
rect 4408 10310 7802 10362
rect 7854 10310 7866 10362
rect 7918 10310 7930 10362
rect 7982 10310 7994 10362
rect 8046 10310 8058 10362
rect 8110 10310 11504 10362
rect 11556 10310 11568 10362
rect 11620 10310 11632 10362
rect 11684 10310 11696 10362
rect 11748 10310 11760 10362
rect 11812 10310 15206 10362
rect 15258 10310 15270 10362
rect 15322 10310 15334 10362
rect 15386 10310 15398 10362
rect 15450 10310 15462 10362
rect 15514 10310 15520 10362
rect 552 10288 15520 10310
rect 6270 10208 6276 10260
rect 6328 10208 6334 10260
rect 10226 10208 10232 10260
rect 10284 10208 10290 10260
rect 8202 10140 8208 10192
rect 8260 10140 8266 10192
rect 8754 10072 8760 10124
rect 8812 10072 8818 10124
rect 9122 10072 9128 10124
rect 9180 10072 9186 10124
rect 10318 10072 10324 10124
rect 10376 10072 10382 10124
rect 6914 10004 6920 10056
rect 6972 10004 6978 10056
rect 7374 9868 7380 9920
rect 7432 9868 7438 9920
rect 552 9818 15364 9840
rect 552 9766 2249 9818
rect 2301 9766 2313 9818
rect 2365 9766 2377 9818
rect 2429 9766 2441 9818
rect 2493 9766 2505 9818
rect 2557 9766 5951 9818
rect 6003 9766 6015 9818
rect 6067 9766 6079 9818
rect 6131 9766 6143 9818
rect 6195 9766 6207 9818
rect 6259 9766 9653 9818
rect 9705 9766 9717 9818
rect 9769 9766 9781 9818
rect 9833 9766 9845 9818
rect 9897 9766 9909 9818
rect 9961 9766 13355 9818
rect 13407 9766 13419 9818
rect 13471 9766 13483 9818
rect 13535 9766 13547 9818
rect 13599 9766 13611 9818
rect 13663 9766 15364 9818
rect 552 9744 15364 9766
rect 6273 9639 6331 9645
rect 6273 9605 6285 9639
rect 6319 9636 6331 9639
rect 6914 9636 6920 9648
rect 6319 9608 6920 9636
rect 6319 9605 6331 9608
rect 6273 9599 6331 9605
rect 6914 9596 6920 9608
rect 6972 9596 6978 9648
rect 8386 9568 8392 9580
rect 6472 9540 8392 9568
rect 6472 9509 6500 9540
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 6457 9503 6515 9509
rect 6457 9469 6469 9503
rect 6503 9469 6515 9503
rect 6457 9463 6515 9469
rect 6638 9460 6644 9512
rect 6696 9460 6702 9512
rect 6733 9503 6791 9509
rect 6733 9469 6745 9503
rect 6779 9500 6791 9503
rect 7374 9500 7380 9512
rect 6779 9472 7380 9500
rect 6779 9469 6791 9472
rect 6733 9463 6791 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 552 9274 15520 9296
rect 552 9222 4100 9274
rect 4152 9222 4164 9274
rect 4216 9222 4228 9274
rect 4280 9222 4292 9274
rect 4344 9222 4356 9274
rect 4408 9222 7802 9274
rect 7854 9222 7866 9274
rect 7918 9222 7930 9274
rect 7982 9222 7994 9274
rect 8046 9222 8058 9274
rect 8110 9222 11504 9274
rect 11556 9222 11568 9274
rect 11620 9222 11632 9274
rect 11684 9222 11696 9274
rect 11748 9222 11760 9274
rect 11812 9222 15206 9274
rect 15258 9222 15270 9274
rect 15322 9222 15334 9274
rect 15386 9222 15398 9274
rect 15450 9222 15462 9274
rect 15514 9222 15520 9274
rect 552 9200 15520 9222
rect 552 8730 15364 8752
rect 552 8678 2249 8730
rect 2301 8678 2313 8730
rect 2365 8678 2377 8730
rect 2429 8678 2441 8730
rect 2493 8678 2505 8730
rect 2557 8678 5951 8730
rect 6003 8678 6015 8730
rect 6067 8678 6079 8730
rect 6131 8678 6143 8730
rect 6195 8678 6207 8730
rect 6259 8678 9653 8730
rect 9705 8678 9717 8730
rect 9769 8678 9781 8730
rect 9833 8678 9845 8730
rect 9897 8678 9909 8730
rect 9961 8678 13355 8730
rect 13407 8678 13419 8730
rect 13471 8678 13483 8730
rect 13535 8678 13547 8730
rect 13599 8678 13611 8730
rect 13663 8678 15364 8730
rect 552 8656 15364 8678
rect 552 8186 15520 8208
rect 552 8134 4100 8186
rect 4152 8134 4164 8186
rect 4216 8134 4228 8186
rect 4280 8134 4292 8186
rect 4344 8134 4356 8186
rect 4408 8134 7802 8186
rect 7854 8134 7866 8186
rect 7918 8134 7930 8186
rect 7982 8134 7994 8186
rect 8046 8134 8058 8186
rect 8110 8134 11504 8186
rect 11556 8134 11568 8186
rect 11620 8134 11632 8186
rect 11684 8134 11696 8186
rect 11748 8134 11760 8186
rect 11812 8134 15206 8186
rect 15258 8134 15270 8186
rect 15322 8134 15334 8186
rect 15386 8134 15398 8186
rect 15450 8134 15462 8186
rect 15514 8134 15520 8186
rect 552 8112 15520 8134
rect 552 7642 15364 7664
rect 552 7590 2249 7642
rect 2301 7590 2313 7642
rect 2365 7590 2377 7642
rect 2429 7590 2441 7642
rect 2493 7590 2505 7642
rect 2557 7590 5951 7642
rect 6003 7590 6015 7642
rect 6067 7590 6079 7642
rect 6131 7590 6143 7642
rect 6195 7590 6207 7642
rect 6259 7590 9653 7642
rect 9705 7590 9717 7642
rect 9769 7590 9781 7642
rect 9833 7590 9845 7642
rect 9897 7590 9909 7642
rect 9961 7590 13355 7642
rect 13407 7590 13419 7642
rect 13471 7590 13483 7642
rect 13535 7590 13547 7642
rect 13599 7590 13611 7642
rect 13663 7590 15364 7642
rect 552 7568 15364 7590
rect 552 7098 15520 7120
rect 552 7046 4100 7098
rect 4152 7046 4164 7098
rect 4216 7046 4228 7098
rect 4280 7046 4292 7098
rect 4344 7046 4356 7098
rect 4408 7046 7802 7098
rect 7854 7046 7866 7098
rect 7918 7046 7930 7098
rect 7982 7046 7994 7098
rect 8046 7046 8058 7098
rect 8110 7046 11504 7098
rect 11556 7046 11568 7098
rect 11620 7046 11632 7098
rect 11684 7046 11696 7098
rect 11748 7046 11760 7098
rect 11812 7046 15206 7098
rect 15258 7046 15270 7098
rect 15322 7046 15334 7098
rect 15386 7046 15398 7098
rect 15450 7046 15462 7098
rect 15514 7046 15520 7098
rect 552 7024 15520 7046
rect 552 6554 15364 6576
rect 552 6502 2249 6554
rect 2301 6502 2313 6554
rect 2365 6502 2377 6554
rect 2429 6502 2441 6554
rect 2493 6502 2505 6554
rect 2557 6502 5951 6554
rect 6003 6502 6015 6554
rect 6067 6502 6079 6554
rect 6131 6502 6143 6554
rect 6195 6502 6207 6554
rect 6259 6502 9653 6554
rect 9705 6502 9717 6554
rect 9769 6502 9781 6554
rect 9833 6502 9845 6554
rect 9897 6502 9909 6554
rect 9961 6502 13355 6554
rect 13407 6502 13419 6554
rect 13471 6502 13483 6554
rect 13535 6502 13547 6554
rect 13599 6502 13611 6554
rect 13663 6502 15364 6554
rect 552 6480 15364 6502
rect 552 6010 15520 6032
rect 552 5958 4100 6010
rect 4152 5958 4164 6010
rect 4216 5958 4228 6010
rect 4280 5958 4292 6010
rect 4344 5958 4356 6010
rect 4408 5958 7802 6010
rect 7854 5958 7866 6010
rect 7918 5958 7930 6010
rect 7982 5958 7994 6010
rect 8046 5958 8058 6010
rect 8110 5958 11504 6010
rect 11556 5958 11568 6010
rect 11620 5958 11632 6010
rect 11684 5958 11696 6010
rect 11748 5958 11760 6010
rect 11812 5958 15206 6010
rect 15258 5958 15270 6010
rect 15322 5958 15334 6010
rect 15386 5958 15398 6010
rect 15450 5958 15462 6010
rect 15514 5958 15520 6010
rect 552 5936 15520 5958
rect 552 5466 15364 5488
rect 552 5414 2249 5466
rect 2301 5414 2313 5466
rect 2365 5414 2377 5466
rect 2429 5414 2441 5466
rect 2493 5414 2505 5466
rect 2557 5414 5951 5466
rect 6003 5414 6015 5466
rect 6067 5414 6079 5466
rect 6131 5414 6143 5466
rect 6195 5414 6207 5466
rect 6259 5414 9653 5466
rect 9705 5414 9717 5466
rect 9769 5414 9781 5466
rect 9833 5414 9845 5466
rect 9897 5414 9909 5466
rect 9961 5414 13355 5466
rect 13407 5414 13419 5466
rect 13471 5414 13483 5466
rect 13535 5414 13547 5466
rect 13599 5414 13611 5466
rect 13663 5414 15364 5466
rect 552 5392 15364 5414
rect 552 4922 15520 4944
rect 552 4870 4100 4922
rect 4152 4870 4164 4922
rect 4216 4870 4228 4922
rect 4280 4870 4292 4922
rect 4344 4870 4356 4922
rect 4408 4870 7802 4922
rect 7854 4870 7866 4922
rect 7918 4870 7930 4922
rect 7982 4870 7994 4922
rect 8046 4870 8058 4922
rect 8110 4870 11504 4922
rect 11556 4870 11568 4922
rect 11620 4870 11632 4922
rect 11684 4870 11696 4922
rect 11748 4870 11760 4922
rect 11812 4870 15206 4922
rect 15258 4870 15270 4922
rect 15322 4870 15334 4922
rect 15386 4870 15398 4922
rect 15450 4870 15462 4922
rect 15514 4870 15520 4922
rect 552 4848 15520 4870
rect 552 4378 15364 4400
rect 552 4326 2249 4378
rect 2301 4326 2313 4378
rect 2365 4326 2377 4378
rect 2429 4326 2441 4378
rect 2493 4326 2505 4378
rect 2557 4326 5951 4378
rect 6003 4326 6015 4378
rect 6067 4326 6079 4378
rect 6131 4326 6143 4378
rect 6195 4326 6207 4378
rect 6259 4326 9653 4378
rect 9705 4326 9717 4378
rect 9769 4326 9781 4378
rect 9833 4326 9845 4378
rect 9897 4326 9909 4378
rect 9961 4326 13355 4378
rect 13407 4326 13419 4378
rect 13471 4326 13483 4378
rect 13535 4326 13547 4378
rect 13599 4326 13611 4378
rect 13663 4326 15364 4378
rect 552 4304 15364 4326
rect 552 3834 15520 3856
rect 552 3782 4100 3834
rect 4152 3782 4164 3834
rect 4216 3782 4228 3834
rect 4280 3782 4292 3834
rect 4344 3782 4356 3834
rect 4408 3782 7802 3834
rect 7854 3782 7866 3834
rect 7918 3782 7930 3834
rect 7982 3782 7994 3834
rect 8046 3782 8058 3834
rect 8110 3782 11504 3834
rect 11556 3782 11568 3834
rect 11620 3782 11632 3834
rect 11684 3782 11696 3834
rect 11748 3782 11760 3834
rect 11812 3782 15206 3834
rect 15258 3782 15270 3834
rect 15322 3782 15334 3834
rect 15386 3782 15398 3834
rect 15450 3782 15462 3834
rect 15514 3782 15520 3834
rect 552 3760 15520 3782
rect 552 3290 15364 3312
rect 552 3238 2249 3290
rect 2301 3238 2313 3290
rect 2365 3238 2377 3290
rect 2429 3238 2441 3290
rect 2493 3238 2505 3290
rect 2557 3238 5951 3290
rect 6003 3238 6015 3290
rect 6067 3238 6079 3290
rect 6131 3238 6143 3290
rect 6195 3238 6207 3290
rect 6259 3238 9653 3290
rect 9705 3238 9717 3290
rect 9769 3238 9781 3290
rect 9833 3238 9845 3290
rect 9897 3238 9909 3290
rect 9961 3238 13355 3290
rect 13407 3238 13419 3290
rect 13471 3238 13483 3290
rect 13535 3238 13547 3290
rect 13599 3238 13611 3290
rect 13663 3238 15364 3290
rect 552 3216 15364 3238
rect 552 2746 15520 2768
rect 552 2694 4100 2746
rect 4152 2694 4164 2746
rect 4216 2694 4228 2746
rect 4280 2694 4292 2746
rect 4344 2694 4356 2746
rect 4408 2694 7802 2746
rect 7854 2694 7866 2746
rect 7918 2694 7930 2746
rect 7982 2694 7994 2746
rect 8046 2694 8058 2746
rect 8110 2694 11504 2746
rect 11556 2694 11568 2746
rect 11620 2694 11632 2746
rect 11684 2694 11696 2746
rect 11748 2694 11760 2746
rect 11812 2694 15206 2746
rect 15258 2694 15270 2746
rect 15322 2694 15334 2746
rect 15386 2694 15398 2746
rect 15450 2694 15462 2746
rect 15514 2694 15520 2746
rect 552 2672 15520 2694
rect 552 2202 15364 2224
rect 552 2150 2249 2202
rect 2301 2150 2313 2202
rect 2365 2150 2377 2202
rect 2429 2150 2441 2202
rect 2493 2150 2505 2202
rect 2557 2150 5951 2202
rect 6003 2150 6015 2202
rect 6067 2150 6079 2202
rect 6131 2150 6143 2202
rect 6195 2150 6207 2202
rect 6259 2150 9653 2202
rect 9705 2150 9717 2202
rect 9769 2150 9781 2202
rect 9833 2150 9845 2202
rect 9897 2150 9909 2202
rect 9961 2150 13355 2202
rect 13407 2150 13419 2202
rect 13471 2150 13483 2202
rect 13535 2150 13547 2202
rect 13599 2150 13611 2202
rect 13663 2150 15364 2202
rect 552 2128 15364 2150
rect 552 1658 15520 1680
rect 552 1606 4100 1658
rect 4152 1606 4164 1658
rect 4216 1606 4228 1658
rect 4280 1606 4292 1658
rect 4344 1606 4356 1658
rect 4408 1606 7802 1658
rect 7854 1606 7866 1658
rect 7918 1606 7930 1658
rect 7982 1606 7994 1658
rect 8046 1606 8058 1658
rect 8110 1606 11504 1658
rect 11556 1606 11568 1658
rect 11620 1606 11632 1658
rect 11684 1606 11696 1658
rect 11748 1606 11760 1658
rect 11812 1606 15206 1658
rect 15258 1606 15270 1658
rect 15322 1606 15334 1658
rect 15386 1606 15398 1658
rect 15450 1606 15462 1658
rect 15514 1606 15520 1658
rect 552 1584 15520 1606
rect 552 1114 15364 1136
rect 552 1062 2249 1114
rect 2301 1062 2313 1114
rect 2365 1062 2377 1114
rect 2429 1062 2441 1114
rect 2493 1062 2505 1114
rect 2557 1062 5951 1114
rect 6003 1062 6015 1114
rect 6067 1062 6079 1114
rect 6131 1062 6143 1114
rect 6195 1062 6207 1114
rect 6259 1062 9653 1114
rect 9705 1062 9717 1114
rect 9769 1062 9781 1114
rect 9833 1062 9845 1114
rect 9897 1062 9909 1114
rect 9961 1062 13355 1114
rect 13407 1062 13419 1114
rect 13471 1062 13483 1114
rect 13535 1062 13547 1114
rect 13599 1062 13611 1114
rect 13663 1062 15364 1114
rect 552 1040 15364 1062
rect 8570 960 8576 1012
rect 8628 960 8634 1012
rect 8478 688 8484 740
rect 8536 688 8542 740
rect 552 570 15520 592
rect 552 518 4100 570
rect 4152 518 4164 570
rect 4216 518 4228 570
rect 4280 518 4292 570
rect 4344 518 4356 570
rect 4408 518 7802 570
rect 7854 518 7866 570
rect 7918 518 7930 570
rect 7982 518 7994 570
rect 8046 518 8058 570
rect 8110 518 11504 570
rect 11556 518 11568 570
rect 11620 518 11632 570
rect 11684 518 11696 570
rect 11748 518 11760 570
rect 11812 518 15206 570
rect 15258 518 15270 570
rect 15322 518 15334 570
rect 15386 518 15398 570
rect 15450 518 15462 570
rect 15514 518 15520 570
rect 552 496 15520 518
rect 8018 416 8024 468
rect 8076 456 8082 468
rect 8478 456 8484 468
rect 8076 428 8484 456
rect 8076 416 8082 428
rect 8478 416 8484 428
rect 8536 416 8542 468
<< via1 >>
rect 2249 15206 2301 15258
rect 2313 15206 2365 15258
rect 2377 15206 2429 15258
rect 2441 15206 2493 15258
rect 2505 15206 2557 15258
rect 5951 15206 6003 15258
rect 6015 15206 6067 15258
rect 6079 15206 6131 15258
rect 6143 15206 6195 15258
rect 6207 15206 6259 15258
rect 9653 15206 9705 15258
rect 9717 15206 9769 15258
rect 9781 15206 9833 15258
rect 9845 15206 9897 15258
rect 9909 15206 9961 15258
rect 13355 15206 13407 15258
rect 13419 15206 13471 15258
rect 13483 15206 13535 15258
rect 13547 15206 13599 15258
rect 13611 15206 13663 15258
rect 8760 15104 8812 15156
rect 1032 14943 1084 14952
rect 1032 14909 1041 14943
rect 1041 14909 1075 14943
rect 1075 14909 1084 14943
rect 1032 14900 1084 14909
rect 8484 14943 8536 14952
rect 8484 14909 8493 14943
rect 8493 14909 8527 14943
rect 8527 14909 8536 14943
rect 8484 14900 8536 14909
rect 3884 14764 3936 14816
rect 4620 14764 4672 14816
rect 4100 14662 4152 14714
rect 4164 14662 4216 14714
rect 4228 14662 4280 14714
rect 4292 14662 4344 14714
rect 4356 14662 4408 14714
rect 7802 14662 7854 14714
rect 7866 14662 7918 14714
rect 7930 14662 7982 14714
rect 7994 14662 8046 14714
rect 8058 14662 8110 14714
rect 11504 14662 11556 14714
rect 11568 14662 11620 14714
rect 11632 14662 11684 14714
rect 11696 14662 11748 14714
rect 11760 14662 11812 14714
rect 15206 14662 15258 14714
rect 15270 14662 15322 14714
rect 15334 14662 15386 14714
rect 15398 14662 15450 14714
rect 15462 14662 15514 14714
rect 4436 14560 4488 14612
rect 5632 14560 5684 14612
rect 7196 14560 7248 14612
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 5816 14424 5868 14476
rect 7104 14492 7156 14544
rect 7748 14492 7800 14544
rect 6276 14467 6328 14476
rect 6276 14433 6285 14467
rect 6285 14433 6319 14467
rect 6319 14433 6328 14467
rect 6276 14424 6328 14433
rect 6368 14424 6420 14476
rect 11796 14492 11848 14544
rect 10784 14467 10836 14476
rect 4896 14356 4948 14408
rect 7012 14399 7064 14408
rect 7012 14365 7021 14399
rect 7021 14365 7055 14399
rect 7055 14365 7064 14399
rect 7012 14356 7064 14365
rect 9036 14399 9088 14408
rect 9036 14365 9045 14399
rect 9045 14365 9079 14399
rect 9079 14365 9088 14399
rect 9036 14356 9088 14365
rect 8208 14288 8260 14340
rect 5632 14220 5684 14272
rect 8484 14263 8536 14272
rect 8484 14229 8493 14263
rect 8493 14229 8527 14263
rect 8527 14229 8536 14263
rect 8484 14220 8536 14229
rect 10784 14433 10793 14467
rect 10793 14433 10827 14467
rect 10827 14433 10836 14467
rect 10784 14424 10836 14433
rect 10968 14467 11020 14476
rect 10968 14433 10977 14467
rect 10977 14433 11011 14467
rect 11011 14433 11020 14467
rect 10968 14424 11020 14433
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 12348 14220 12400 14272
rect 2249 14118 2301 14170
rect 2313 14118 2365 14170
rect 2377 14118 2429 14170
rect 2441 14118 2493 14170
rect 2505 14118 2557 14170
rect 5951 14118 6003 14170
rect 6015 14118 6067 14170
rect 6079 14118 6131 14170
rect 6143 14118 6195 14170
rect 6207 14118 6259 14170
rect 9653 14118 9705 14170
rect 9717 14118 9769 14170
rect 9781 14118 9833 14170
rect 9845 14118 9897 14170
rect 9909 14118 9961 14170
rect 13355 14118 13407 14170
rect 13419 14118 13471 14170
rect 13483 14118 13535 14170
rect 13547 14118 13599 14170
rect 13611 14118 13663 14170
rect 4896 13880 4948 13932
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 7104 14016 7156 14068
rect 6552 13948 6604 14000
rect 7748 14016 7800 14068
rect 10324 14016 10376 14068
rect 11796 14059 11848 14068
rect 11796 14025 11805 14059
rect 11805 14025 11839 14059
rect 11839 14025 11848 14059
rect 11796 14016 11848 14025
rect 8208 13948 8260 14000
rect 10692 13948 10744 14000
rect 8484 13880 8536 13932
rect 12348 13880 12400 13932
rect 5632 13744 5684 13796
rect 6184 13744 6236 13796
rect 8208 13812 8260 13864
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 5540 13676 5592 13728
rect 6920 13676 6972 13728
rect 9220 13744 9272 13796
rect 9864 13744 9916 13796
rect 10784 13812 10836 13864
rect 7656 13676 7708 13728
rect 8484 13676 8536 13728
rect 11336 13676 11388 13728
rect 4100 13574 4152 13626
rect 4164 13574 4216 13626
rect 4228 13574 4280 13626
rect 4292 13574 4344 13626
rect 4356 13574 4408 13626
rect 7802 13574 7854 13626
rect 7866 13574 7918 13626
rect 7930 13574 7982 13626
rect 7994 13574 8046 13626
rect 8058 13574 8110 13626
rect 11504 13574 11556 13626
rect 11568 13574 11620 13626
rect 11632 13574 11684 13626
rect 11696 13574 11748 13626
rect 11760 13574 11812 13626
rect 15206 13574 15258 13626
rect 15270 13574 15322 13626
rect 15334 13574 15386 13626
rect 15398 13574 15450 13626
rect 15462 13574 15514 13626
rect 6184 13472 6236 13524
rect 7012 13472 7064 13524
rect 5172 13404 5224 13456
rect 3884 13379 3936 13388
rect 3884 13345 3893 13379
rect 3893 13345 3927 13379
rect 3927 13345 3936 13379
rect 3884 13336 3936 13345
rect 3056 13311 3108 13320
rect 3056 13277 3065 13311
rect 3065 13277 3099 13311
rect 3099 13277 3108 13311
rect 3056 13268 3108 13277
rect 4988 13311 5040 13320
rect 4988 13277 4997 13311
rect 4997 13277 5031 13311
rect 5031 13277 5040 13311
rect 4988 13268 5040 13277
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 5540 13379 5592 13388
rect 5540 13345 5549 13379
rect 5549 13345 5583 13379
rect 5583 13345 5592 13379
rect 5540 13336 5592 13345
rect 5724 13268 5776 13320
rect 5816 13268 5868 13320
rect 6736 13336 6788 13388
rect 7196 13336 7248 13388
rect 7656 13379 7708 13388
rect 7656 13345 7665 13379
rect 7665 13345 7699 13379
rect 7699 13345 7708 13379
rect 7656 13336 7708 13345
rect 3792 13175 3844 13184
rect 3792 13141 3801 13175
rect 3801 13141 3835 13175
rect 3835 13141 3844 13175
rect 3792 13132 3844 13141
rect 4804 13132 4856 13184
rect 6460 13200 6512 13252
rect 6552 13200 6604 13252
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 7564 13311 7616 13320
rect 7564 13277 7573 13311
rect 7573 13277 7607 13311
rect 7607 13277 7616 13311
rect 9036 13472 9088 13524
rect 10140 13472 10192 13524
rect 11244 13472 11296 13524
rect 8576 13379 8628 13388
rect 8576 13345 8585 13379
rect 8585 13345 8619 13379
rect 8619 13345 8628 13379
rect 8576 13336 8628 13345
rect 7564 13268 7616 13277
rect 8392 13268 8444 13320
rect 9128 13336 9180 13388
rect 9312 13311 9364 13320
rect 9312 13277 9321 13311
rect 9321 13277 9355 13311
rect 9355 13277 9364 13311
rect 9312 13268 9364 13277
rect 9956 13336 10008 13388
rect 10048 13336 10100 13388
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 10692 13379 10744 13388
rect 10692 13345 10701 13379
rect 10701 13345 10735 13379
rect 10735 13345 10744 13379
rect 10692 13336 10744 13345
rect 10784 13336 10836 13388
rect 10324 13268 10376 13320
rect 5172 13132 5224 13184
rect 6644 13175 6696 13184
rect 6644 13141 6653 13175
rect 6653 13141 6687 13175
rect 6687 13141 6696 13175
rect 6644 13132 6696 13141
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 7472 13243 7524 13252
rect 7472 13209 7481 13243
rect 7481 13209 7515 13243
rect 7515 13209 7524 13243
rect 7472 13200 7524 13209
rect 9864 13200 9916 13252
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 7656 13132 7708 13184
rect 8208 13132 8260 13184
rect 9220 13132 9272 13184
rect 9956 13132 10008 13184
rect 10232 13175 10284 13184
rect 10232 13141 10241 13175
rect 10241 13141 10275 13175
rect 10275 13141 10284 13175
rect 10232 13132 10284 13141
rect 10692 13132 10744 13184
rect 2249 13030 2301 13082
rect 2313 13030 2365 13082
rect 2377 13030 2429 13082
rect 2441 13030 2493 13082
rect 2505 13030 2557 13082
rect 5951 13030 6003 13082
rect 6015 13030 6067 13082
rect 6079 13030 6131 13082
rect 6143 13030 6195 13082
rect 6207 13030 6259 13082
rect 9653 13030 9705 13082
rect 9717 13030 9769 13082
rect 9781 13030 9833 13082
rect 9845 13030 9897 13082
rect 9909 13030 9961 13082
rect 13355 13030 13407 13082
rect 13419 13030 13471 13082
rect 13483 13030 13535 13082
rect 13547 13030 13599 13082
rect 13611 13030 13663 13082
rect 4896 12928 4948 12980
rect 4988 12928 5040 12980
rect 6092 12928 6144 12980
rect 7012 12928 7064 12980
rect 8760 12928 8812 12980
rect 10416 12928 10468 12980
rect 10784 12928 10836 12980
rect 13084 12928 13136 12980
rect 4804 12792 4856 12844
rect 5632 12792 5684 12844
rect 7472 12860 7524 12912
rect 8484 12860 8536 12912
rect 6460 12699 6512 12708
rect 6460 12665 6469 12699
rect 6469 12665 6503 12699
rect 6503 12665 6512 12699
rect 6460 12656 6512 12665
rect 8392 12724 8444 12776
rect 8576 12724 8628 12776
rect 8944 12767 8996 12776
rect 8944 12733 8953 12767
rect 8953 12733 8987 12767
rect 8987 12733 8996 12767
rect 8944 12724 8996 12733
rect 9680 12724 9732 12776
rect 9864 12724 9916 12776
rect 12716 12767 12768 12776
rect 12716 12733 12725 12767
rect 12725 12733 12759 12767
rect 12759 12733 12768 12767
rect 12716 12724 12768 12733
rect 8208 12699 8260 12708
rect 8208 12665 8217 12699
rect 8217 12665 8251 12699
rect 8251 12665 8260 12699
rect 8208 12656 8260 12665
rect 6092 12588 6144 12640
rect 10140 12656 10192 12708
rect 4100 12486 4152 12538
rect 4164 12486 4216 12538
rect 4228 12486 4280 12538
rect 4292 12486 4344 12538
rect 4356 12486 4408 12538
rect 7802 12486 7854 12538
rect 7866 12486 7918 12538
rect 7930 12486 7982 12538
rect 7994 12486 8046 12538
rect 8058 12486 8110 12538
rect 11504 12486 11556 12538
rect 11568 12486 11620 12538
rect 11632 12486 11684 12538
rect 11696 12486 11748 12538
rect 11760 12486 11812 12538
rect 15206 12486 15258 12538
rect 15270 12486 15322 12538
rect 15334 12486 15386 12538
rect 15398 12486 15450 12538
rect 15462 12486 15514 12538
rect 3792 12316 3844 12368
rect 4896 12384 4948 12436
rect 5816 12384 5868 12436
rect 6736 12427 6788 12436
rect 4436 12316 4488 12368
rect 4712 12316 4764 12368
rect 5724 12316 5776 12368
rect 5816 12248 5868 12300
rect 6736 12393 6745 12427
rect 6745 12393 6779 12427
rect 6779 12393 6788 12427
rect 6736 12384 6788 12393
rect 7656 12384 7708 12436
rect 6552 12316 6604 12368
rect 6092 12291 6144 12300
rect 6092 12257 6101 12291
rect 6101 12257 6135 12291
rect 6135 12257 6144 12291
rect 6092 12248 6144 12257
rect 6644 12248 6696 12300
rect 3056 12180 3108 12232
rect 6552 12180 6604 12232
rect 6368 12112 6420 12164
rect 6920 12291 6972 12300
rect 6920 12257 6929 12291
rect 6929 12257 6963 12291
rect 6963 12257 6972 12291
rect 6920 12248 6972 12257
rect 8208 12248 8260 12300
rect 8484 12384 8536 12436
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 8576 12316 8628 12368
rect 9312 12316 9364 12368
rect 7564 12180 7616 12232
rect 8944 12248 8996 12300
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 10416 12359 10468 12368
rect 10416 12325 10425 12359
rect 10425 12325 10459 12359
rect 10459 12325 10468 12359
rect 10416 12316 10468 12325
rect 9680 12248 9732 12300
rect 10324 12291 10376 12300
rect 10324 12257 10333 12291
rect 10333 12257 10367 12291
rect 10367 12257 10376 12291
rect 10324 12248 10376 12257
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 12624 12248 12676 12300
rect 10048 12223 10100 12232
rect 10048 12189 10057 12223
rect 10057 12189 10091 12223
rect 10091 12189 10100 12223
rect 10048 12180 10100 12189
rect 10968 12223 11020 12232
rect 10968 12189 10977 12223
rect 10977 12189 11011 12223
rect 11011 12189 11020 12223
rect 10968 12180 11020 12189
rect 10508 12112 10560 12164
rect 8208 12044 8260 12096
rect 8392 12044 8444 12096
rect 9312 12087 9364 12096
rect 9312 12053 9321 12087
rect 9321 12053 9355 12087
rect 9355 12053 9364 12087
rect 9312 12044 9364 12053
rect 2249 11942 2301 11994
rect 2313 11942 2365 11994
rect 2377 11942 2429 11994
rect 2441 11942 2493 11994
rect 2505 11942 2557 11994
rect 5951 11942 6003 11994
rect 6015 11942 6067 11994
rect 6079 11942 6131 11994
rect 6143 11942 6195 11994
rect 6207 11942 6259 11994
rect 9653 11942 9705 11994
rect 9717 11942 9769 11994
rect 9781 11942 9833 11994
rect 9845 11942 9897 11994
rect 9909 11942 9961 11994
rect 13355 11942 13407 11994
rect 13419 11942 13471 11994
rect 13483 11942 13535 11994
rect 13547 11942 13599 11994
rect 13611 11942 13663 11994
rect 4712 11883 4764 11892
rect 4712 11849 4721 11883
rect 4721 11849 4755 11883
rect 4755 11849 4764 11883
rect 4712 11840 4764 11849
rect 7564 11840 7616 11892
rect 8300 11840 8352 11892
rect 5816 11772 5868 11824
rect 6368 11772 6420 11824
rect 10048 11840 10100 11892
rect 12624 11883 12676 11892
rect 12624 11849 12633 11883
rect 12633 11849 12667 11883
rect 12667 11849 12676 11883
rect 12624 11840 12676 11849
rect 15016 11840 15068 11892
rect 10232 11772 10284 11824
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 5540 11679 5592 11688
rect 5540 11645 5549 11679
rect 5549 11645 5583 11679
rect 5583 11645 5592 11679
rect 5540 11636 5592 11645
rect 5632 11636 5684 11688
rect 6368 11636 6420 11688
rect 6552 11679 6604 11688
rect 6552 11645 6561 11679
rect 6561 11645 6595 11679
rect 6595 11645 6604 11679
rect 6552 11636 6604 11645
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 6828 11636 6880 11688
rect 7656 11679 7708 11688
rect 7656 11645 7695 11679
rect 7695 11645 7708 11679
rect 7656 11636 7708 11645
rect 13084 11704 13136 11756
rect 9404 11568 9456 11620
rect 9956 11568 10008 11620
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 12532 11679 12584 11688
rect 12532 11645 12541 11679
rect 12541 11645 12575 11679
rect 12575 11645 12584 11679
rect 12532 11636 12584 11645
rect 12716 11636 12768 11688
rect 5356 11543 5408 11552
rect 5356 11509 5365 11543
rect 5365 11509 5399 11543
rect 5399 11509 5408 11543
rect 5356 11500 5408 11509
rect 6920 11500 6972 11552
rect 7380 11500 7432 11552
rect 9128 11500 9180 11552
rect 10508 11500 10560 11552
rect 10968 11500 11020 11552
rect 4100 11398 4152 11450
rect 4164 11398 4216 11450
rect 4228 11398 4280 11450
rect 4292 11398 4344 11450
rect 4356 11398 4408 11450
rect 7802 11398 7854 11450
rect 7866 11398 7918 11450
rect 7930 11398 7982 11450
rect 7994 11398 8046 11450
rect 8058 11398 8110 11450
rect 11504 11398 11556 11450
rect 11568 11398 11620 11450
rect 11632 11398 11684 11450
rect 11696 11398 11748 11450
rect 11760 11398 11812 11450
rect 15206 11398 15258 11450
rect 15270 11398 15322 11450
rect 15334 11398 15386 11450
rect 15398 11398 15450 11450
rect 15462 11398 15514 11450
rect 6276 11296 6328 11348
rect 6828 11296 6880 11348
rect 9036 11296 9088 11348
rect 4160 11228 4212 11280
rect 4436 11228 4488 11280
rect 8668 11228 8720 11280
rect 9312 11228 9364 11280
rect 9864 11228 9916 11280
rect 12164 11296 12216 11348
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 11520 11228 11572 11280
rect 7012 11160 7064 11212
rect 7288 11160 7340 11212
rect 5356 11092 5408 11144
rect 7380 11092 7432 11144
rect 8576 11203 8628 11212
rect 8576 11169 8585 11203
rect 8585 11169 8619 11203
rect 8619 11169 8628 11203
rect 8576 11160 8628 11169
rect 9036 11203 9088 11212
rect 9036 11169 9045 11203
rect 9045 11169 9079 11203
rect 9079 11169 9088 11203
rect 9036 11160 9088 11169
rect 9128 11203 9180 11212
rect 9128 11169 9137 11203
rect 9137 11169 9171 11203
rect 9171 11169 9180 11203
rect 9128 11160 9180 11169
rect 9496 11160 9548 11212
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 10232 11203 10284 11212
rect 10232 11169 10241 11203
rect 10241 11169 10275 11203
rect 10275 11169 10284 11203
rect 10232 11160 10284 11169
rect 10508 11160 10560 11212
rect 8484 11092 8536 11144
rect 6920 11024 6972 11076
rect 10048 11092 10100 11144
rect 10968 11135 11020 11144
rect 10968 11101 10977 11135
rect 10977 11101 11011 11135
rect 11011 11101 11020 11135
rect 10968 11092 11020 11101
rect 8760 10999 8812 11008
rect 8760 10965 8769 10999
rect 8769 10965 8803 10999
rect 8803 10965 8812 10999
rect 8760 10956 8812 10965
rect 9220 10999 9272 11008
rect 9220 10965 9229 10999
rect 9229 10965 9263 10999
rect 9263 10965 9272 10999
rect 9220 10956 9272 10965
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 9864 10999 9916 11008
rect 9864 10965 9873 10999
rect 9873 10965 9907 10999
rect 9907 10965 9916 10999
rect 9864 10956 9916 10965
rect 2249 10854 2301 10906
rect 2313 10854 2365 10906
rect 2377 10854 2429 10906
rect 2441 10854 2493 10906
rect 2505 10854 2557 10906
rect 5951 10854 6003 10906
rect 6015 10854 6067 10906
rect 6079 10854 6131 10906
rect 6143 10854 6195 10906
rect 6207 10854 6259 10906
rect 9653 10854 9705 10906
rect 9717 10854 9769 10906
rect 9781 10854 9833 10906
rect 9845 10854 9897 10906
rect 9909 10854 9961 10906
rect 13355 10854 13407 10906
rect 13419 10854 13471 10906
rect 13483 10854 13535 10906
rect 13547 10854 13599 10906
rect 13611 10854 13663 10906
rect 4160 10616 4212 10668
rect 7656 10616 7708 10668
rect 9496 10752 9548 10804
rect 10048 10752 10100 10804
rect 10324 10752 10376 10804
rect 11520 10795 11572 10804
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 10968 10616 11020 10668
rect 6276 10548 6328 10600
rect 7012 10548 7064 10600
rect 6920 10480 6972 10532
rect 8208 10412 8260 10464
rect 8392 10455 8444 10464
rect 8392 10421 8401 10455
rect 8401 10421 8435 10455
rect 8435 10421 8444 10455
rect 8392 10412 8444 10421
rect 9128 10591 9180 10600
rect 9128 10557 9137 10591
rect 9137 10557 9171 10591
rect 9171 10557 9180 10591
rect 9128 10548 9180 10557
rect 9220 10548 9272 10600
rect 10324 10548 10376 10600
rect 12532 10548 12584 10600
rect 10232 10480 10284 10532
rect 10324 10412 10376 10464
rect 4100 10310 4152 10362
rect 4164 10310 4216 10362
rect 4228 10310 4280 10362
rect 4292 10310 4344 10362
rect 4356 10310 4408 10362
rect 7802 10310 7854 10362
rect 7866 10310 7918 10362
rect 7930 10310 7982 10362
rect 7994 10310 8046 10362
rect 8058 10310 8110 10362
rect 11504 10310 11556 10362
rect 11568 10310 11620 10362
rect 11632 10310 11684 10362
rect 11696 10310 11748 10362
rect 11760 10310 11812 10362
rect 15206 10310 15258 10362
rect 15270 10310 15322 10362
rect 15334 10310 15386 10362
rect 15398 10310 15450 10362
rect 15462 10310 15514 10362
rect 6276 10251 6328 10260
rect 6276 10217 6285 10251
rect 6285 10217 6319 10251
rect 6319 10217 6328 10251
rect 6276 10208 6328 10217
rect 10232 10251 10284 10260
rect 10232 10217 10241 10251
rect 10241 10217 10275 10251
rect 10275 10217 10284 10251
rect 10232 10208 10284 10217
rect 8208 10140 8260 10192
rect 8760 10115 8812 10124
rect 8760 10081 8769 10115
rect 8769 10081 8803 10115
rect 8803 10081 8812 10115
rect 8760 10072 8812 10081
rect 9128 10115 9180 10124
rect 9128 10081 9137 10115
rect 9137 10081 9171 10115
rect 9171 10081 9180 10115
rect 9128 10072 9180 10081
rect 10324 10115 10376 10124
rect 10324 10081 10333 10115
rect 10333 10081 10367 10115
rect 10367 10081 10376 10115
rect 10324 10072 10376 10081
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 7380 9911 7432 9920
rect 7380 9877 7389 9911
rect 7389 9877 7423 9911
rect 7423 9877 7432 9911
rect 7380 9868 7432 9877
rect 2249 9766 2301 9818
rect 2313 9766 2365 9818
rect 2377 9766 2429 9818
rect 2441 9766 2493 9818
rect 2505 9766 2557 9818
rect 5951 9766 6003 9818
rect 6015 9766 6067 9818
rect 6079 9766 6131 9818
rect 6143 9766 6195 9818
rect 6207 9766 6259 9818
rect 9653 9766 9705 9818
rect 9717 9766 9769 9818
rect 9781 9766 9833 9818
rect 9845 9766 9897 9818
rect 9909 9766 9961 9818
rect 13355 9766 13407 9818
rect 13419 9766 13471 9818
rect 13483 9766 13535 9818
rect 13547 9766 13599 9818
rect 13611 9766 13663 9818
rect 6920 9596 6972 9648
rect 8392 9528 8444 9580
rect 6644 9503 6696 9512
rect 6644 9469 6653 9503
rect 6653 9469 6687 9503
rect 6687 9469 6696 9503
rect 6644 9460 6696 9469
rect 7380 9460 7432 9512
rect 4100 9222 4152 9274
rect 4164 9222 4216 9274
rect 4228 9222 4280 9274
rect 4292 9222 4344 9274
rect 4356 9222 4408 9274
rect 7802 9222 7854 9274
rect 7866 9222 7918 9274
rect 7930 9222 7982 9274
rect 7994 9222 8046 9274
rect 8058 9222 8110 9274
rect 11504 9222 11556 9274
rect 11568 9222 11620 9274
rect 11632 9222 11684 9274
rect 11696 9222 11748 9274
rect 11760 9222 11812 9274
rect 15206 9222 15258 9274
rect 15270 9222 15322 9274
rect 15334 9222 15386 9274
rect 15398 9222 15450 9274
rect 15462 9222 15514 9274
rect 2249 8678 2301 8730
rect 2313 8678 2365 8730
rect 2377 8678 2429 8730
rect 2441 8678 2493 8730
rect 2505 8678 2557 8730
rect 5951 8678 6003 8730
rect 6015 8678 6067 8730
rect 6079 8678 6131 8730
rect 6143 8678 6195 8730
rect 6207 8678 6259 8730
rect 9653 8678 9705 8730
rect 9717 8678 9769 8730
rect 9781 8678 9833 8730
rect 9845 8678 9897 8730
rect 9909 8678 9961 8730
rect 13355 8678 13407 8730
rect 13419 8678 13471 8730
rect 13483 8678 13535 8730
rect 13547 8678 13599 8730
rect 13611 8678 13663 8730
rect 4100 8134 4152 8186
rect 4164 8134 4216 8186
rect 4228 8134 4280 8186
rect 4292 8134 4344 8186
rect 4356 8134 4408 8186
rect 7802 8134 7854 8186
rect 7866 8134 7918 8186
rect 7930 8134 7982 8186
rect 7994 8134 8046 8186
rect 8058 8134 8110 8186
rect 11504 8134 11556 8186
rect 11568 8134 11620 8186
rect 11632 8134 11684 8186
rect 11696 8134 11748 8186
rect 11760 8134 11812 8186
rect 15206 8134 15258 8186
rect 15270 8134 15322 8186
rect 15334 8134 15386 8186
rect 15398 8134 15450 8186
rect 15462 8134 15514 8186
rect 2249 7590 2301 7642
rect 2313 7590 2365 7642
rect 2377 7590 2429 7642
rect 2441 7590 2493 7642
rect 2505 7590 2557 7642
rect 5951 7590 6003 7642
rect 6015 7590 6067 7642
rect 6079 7590 6131 7642
rect 6143 7590 6195 7642
rect 6207 7590 6259 7642
rect 9653 7590 9705 7642
rect 9717 7590 9769 7642
rect 9781 7590 9833 7642
rect 9845 7590 9897 7642
rect 9909 7590 9961 7642
rect 13355 7590 13407 7642
rect 13419 7590 13471 7642
rect 13483 7590 13535 7642
rect 13547 7590 13599 7642
rect 13611 7590 13663 7642
rect 4100 7046 4152 7098
rect 4164 7046 4216 7098
rect 4228 7046 4280 7098
rect 4292 7046 4344 7098
rect 4356 7046 4408 7098
rect 7802 7046 7854 7098
rect 7866 7046 7918 7098
rect 7930 7046 7982 7098
rect 7994 7046 8046 7098
rect 8058 7046 8110 7098
rect 11504 7046 11556 7098
rect 11568 7046 11620 7098
rect 11632 7046 11684 7098
rect 11696 7046 11748 7098
rect 11760 7046 11812 7098
rect 15206 7046 15258 7098
rect 15270 7046 15322 7098
rect 15334 7046 15386 7098
rect 15398 7046 15450 7098
rect 15462 7046 15514 7098
rect 2249 6502 2301 6554
rect 2313 6502 2365 6554
rect 2377 6502 2429 6554
rect 2441 6502 2493 6554
rect 2505 6502 2557 6554
rect 5951 6502 6003 6554
rect 6015 6502 6067 6554
rect 6079 6502 6131 6554
rect 6143 6502 6195 6554
rect 6207 6502 6259 6554
rect 9653 6502 9705 6554
rect 9717 6502 9769 6554
rect 9781 6502 9833 6554
rect 9845 6502 9897 6554
rect 9909 6502 9961 6554
rect 13355 6502 13407 6554
rect 13419 6502 13471 6554
rect 13483 6502 13535 6554
rect 13547 6502 13599 6554
rect 13611 6502 13663 6554
rect 4100 5958 4152 6010
rect 4164 5958 4216 6010
rect 4228 5958 4280 6010
rect 4292 5958 4344 6010
rect 4356 5958 4408 6010
rect 7802 5958 7854 6010
rect 7866 5958 7918 6010
rect 7930 5958 7982 6010
rect 7994 5958 8046 6010
rect 8058 5958 8110 6010
rect 11504 5958 11556 6010
rect 11568 5958 11620 6010
rect 11632 5958 11684 6010
rect 11696 5958 11748 6010
rect 11760 5958 11812 6010
rect 15206 5958 15258 6010
rect 15270 5958 15322 6010
rect 15334 5958 15386 6010
rect 15398 5958 15450 6010
rect 15462 5958 15514 6010
rect 2249 5414 2301 5466
rect 2313 5414 2365 5466
rect 2377 5414 2429 5466
rect 2441 5414 2493 5466
rect 2505 5414 2557 5466
rect 5951 5414 6003 5466
rect 6015 5414 6067 5466
rect 6079 5414 6131 5466
rect 6143 5414 6195 5466
rect 6207 5414 6259 5466
rect 9653 5414 9705 5466
rect 9717 5414 9769 5466
rect 9781 5414 9833 5466
rect 9845 5414 9897 5466
rect 9909 5414 9961 5466
rect 13355 5414 13407 5466
rect 13419 5414 13471 5466
rect 13483 5414 13535 5466
rect 13547 5414 13599 5466
rect 13611 5414 13663 5466
rect 4100 4870 4152 4922
rect 4164 4870 4216 4922
rect 4228 4870 4280 4922
rect 4292 4870 4344 4922
rect 4356 4870 4408 4922
rect 7802 4870 7854 4922
rect 7866 4870 7918 4922
rect 7930 4870 7982 4922
rect 7994 4870 8046 4922
rect 8058 4870 8110 4922
rect 11504 4870 11556 4922
rect 11568 4870 11620 4922
rect 11632 4870 11684 4922
rect 11696 4870 11748 4922
rect 11760 4870 11812 4922
rect 15206 4870 15258 4922
rect 15270 4870 15322 4922
rect 15334 4870 15386 4922
rect 15398 4870 15450 4922
rect 15462 4870 15514 4922
rect 2249 4326 2301 4378
rect 2313 4326 2365 4378
rect 2377 4326 2429 4378
rect 2441 4326 2493 4378
rect 2505 4326 2557 4378
rect 5951 4326 6003 4378
rect 6015 4326 6067 4378
rect 6079 4326 6131 4378
rect 6143 4326 6195 4378
rect 6207 4326 6259 4378
rect 9653 4326 9705 4378
rect 9717 4326 9769 4378
rect 9781 4326 9833 4378
rect 9845 4326 9897 4378
rect 9909 4326 9961 4378
rect 13355 4326 13407 4378
rect 13419 4326 13471 4378
rect 13483 4326 13535 4378
rect 13547 4326 13599 4378
rect 13611 4326 13663 4378
rect 4100 3782 4152 3834
rect 4164 3782 4216 3834
rect 4228 3782 4280 3834
rect 4292 3782 4344 3834
rect 4356 3782 4408 3834
rect 7802 3782 7854 3834
rect 7866 3782 7918 3834
rect 7930 3782 7982 3834
rect 7994 3782 8046 3834
rect 8058 3782 8110 3834
rect 11504 3782 11556 3834
rect 11568 3782 11620 3834
rect 11632 3782 11684 3834
rect 11696 3782 11748 3834
rect 11760 3782 11812 3834
rect 15206 3782 15258 3834
rect 15270 3782 15322 3834
rect 15334 3782 15386 3834
rect 15398 3782 15450 3834
rect 15462 3782 15514 3834
rect 2249 3238 2301 3290
rect 2313 3238 2365 3290
rect 2377 3238 2429 3290
rect 2441 3238 2493 3290
rect 2505 3238 2557 3290
rect 5951 3238 6003 3290
rect 6015 3238 6067 3290
rect 6079 3238 6131 3290
rect 6143 3238 6195 3290
rect 6207 3238 6259 3290
rect 9653 3238 9705 3290
rect 9717 3238 9769 3290
rect 9781 3238 9833 3290
rect 9845 3238 9897 3290
rect 9909 3238 9961 3290
rect 13355 3238 13407 3290
rect 13419 3238 13471 3290
rect 13483 3238 13535 3290
rect 13547 3238 13599 3290
rect 13611 3238 13663 3290
rect 4100 2694 4152 2746
rect 4164 2694 4216 2746
rect 4228 2694 4280 2746
rect 4292 2694 4344 2746
rect 4356 2694 4408 2746
rect 7802 2694 7854 2746
rect 7866 2694 7918 2746
rect 7930 2694 7982 2746
rect 7994 2694 8046 2746
rect 8058 2694 8110 2746
rect 11504 2694 11556 2746
rect 11568 2694 11620 2746
rect 11632 2694 11684 2746
rect 11696 2694 11748 2746
rect 11760 2694 11812 2746
rect 15206 2694 15258 2746
rect 15270 2694 15322 2746
rect 15334 2694 15386 2746
rect 15398 2694 15450 2746
rect 15462 2694 15514 2746
rect 2249 2150 2301 2202
rect 2313 2150 2365 2202
rect 2377 2150 2429 2202
rect 2441 2150 2493 2202
rect 2505 2150 2557 2202
rect 5951 2150 6003 2202
rect 6015 2150 6067 2202
rect 6079 2150 6131 2202
rect 6143 2150 6195 2202
rect 6207 2150 6259 2202
rect 9653 2150 9705 2202
rect 9717 2150 9769 2202
rect 9781 2150 9833 2202
rect 9845 2150 9897 2202
rect 9909 2150 9961 2202
rect 13355 2150 13407 2202
rect 13419 2150 13471 2202
rect 13483 2150 13535 2202
rect 13547 2150 13599 2202
rect 13611 2150 13663 2202
rect 4100 1606 4152 1658
rect 4164 1606 4216 1658
rect 4228 1606 4280 1658
rect 4292 1606 4344 1658
rect 4356 1606 4408 1658
rect 7802 1606 7854 1658
rect 7866 1606 7918 1658
rect 7930 1606 7982 1658
rect 7994 1606 8046 1658
rect 8058 1606 8110 1658
rect 11504 1606 11556 1658
rect 11568 1606 11620 1658
rect 11632 1606 11684 1658
rect 11696 1606 11748 1658
rect 11760 1606 11812 1658
rect 15206 1606 15258 1658
rect 15270 1606 15322 1658
rect 15334 1606 15386 1658
rect 15398 1606 15450 1658
rect 15462 1606 15514 1658
rect 2249 1062 2301 1114
rect 2313 1062 2365 1114
rect 2377 1062 2429 1114
rect 2441 1062 2493 1114
rect 2505 1062 2557 1114
rect 5951 1062 6003 1114
rect 6015 1062 6067 1114
rect 6079 1062 6131 1114
rect 6143 1062 6195 1114
rect 6207 1062 6259 1114
rect 9653 1062 9705 1114
rect 9717 1062 9769 1114
rect 9781 1062 9833 1114
rect 9845 1062 9897 1114
rect 9909 1062 9961 1114
rect 13355 1062 13407 1114
rect 13419 1062 13471 1114
rect 13483 1062 13535 1114
rect 13547 1062 13599 1114
rect 13611 1062 13663 1114
rect 8576 1003 8628 1012
rect 8576 969 8585 1003
rect 8585 969 8619 1003
rect 8619 969 8628 1003
rect 8576 960 8628 969
rect 8484 731 8536 740
rect 8484 697 8493 731
rect 8493 697 8527 731
rect 8527 697 8536 731
rect 8484 688 8536 697
rect 4100 518 4152 570
rect 4164 518 4216 570
rect 4228 518 4280 570
rect 4292 518 4344 570
rect 4356 518 4408 570
rect 7802 518 7854 570
rect 7866 518 7918 570
rect 7930 518 7982 570
rect 7994 518 8046 570
rect 8058 518 8110 570
rect 11504 518 11556 570
rect 11568 518 11620 570
rect 11632 518 11684 570
rect 11696 518 11748 570
rect 11760 518 11812 570
rect 15206 518 15258 570
rect 15270 518 15322 570
rect 15334 518 15386 570
rect 15398 518 15450 570
rect 15462 518 15514 570
rect 8024 416 8076 468
rect 8484 416 8536 468
<< metal2 >>
rect 938 15722 994 16000
rect 2502 15722 2558 16000
rect 4066 15722 4122 16000
rect 938 15694 1072 15722
rect 938 15600 994 15694
rect 1044 14958 1072 15694
rect 2502 15694 2728 15722
rect 2502 15600 2558 15694
rect 2249 15260 2557 15269
rect 2249 15258 2255 15260
rect 2311 15258 2335 15260
rect 2391 15258 2415 15260
rect 2471 15258 2495 15260
rect 2551 15258 2557 15260
rect 2311 15206 2313 15258
rect 2493 15206 2495 15258
rect 2249 15204 2255 15206
rect 2311 15204 2335 15206
rect 2391 15204 2415 15206
rect 2471 15204 2495 15206
rect 2551 15204 2557 15206
rect 2249 15195 2557 15204
rect 1032 14952 1084 14958
rect 1032 14894 1084 14900
rect 2249 14172 2557 14181
rect 2249 14170 2255 14172
rect 2311 14170 2335 14172
rect 2391 14170 2415 14172
rect 2471 14170 2495 14172
rect 2551 14170 2557 14172
rect 2311 14118 2313 14170
rect 2493 14118 2495 14170
rect 2249 14116 2255 14118
rect 2311 14116 2335 14118
rect 2391 14116 2415 14118
rect 2471 14116 2495 14118
rect 2551 14116 2557 14118
rect 2249 14107 2557 14116
rect 2249 13084 2557 13093
rect 2249 13082 2255 13084
rect 2311 13082 2335 13084
rect 2391 13082 2415 13084
rect 2471 13082 2495 13084
rect 2551 13082 2557 13084
rect 2311 13030 2313 13082
rect 2493 13030 2495 13082
rect 2249 13028 2255 13030
rect 2311 13028 2335 13030
rect 2391 13028 2415 13030
rect 2471 13028 2495 13030
rect 2551 13028 2557 13030
rect 2249 13019 2557 13028
rect 2700 12345 2728 15694
rect 4066 15694 4476 15722
rect 4066 15600 4122 15694
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 13394 3924 14758
rect 4100 14716 4408 14725
rect 4100 14714 4106 14716
rect 4162 14714 4186 14716
rect 4242 14714 4266 14716
rect 4322 14714 4346 14716
rect 4402 14714 4408 14716
rect 4162 14662 4164 14714
rect 4344 14662 4346 14714
rect 4100 14660 4106 14662
rect 4162 14660 4186 14662
rect 4242 14660 4266 14662
rect 4322 14660 4346 14662
rect 4402 14660 4408 14662
rect 4100 14651 4408 14660
rect 4448 14618 4476 15694
rect 5630 15600 5686 16000
rect 7194 15600 7250 16000
rect 8758 15600 8814 16000
rect 10322 15600 10378 16000
rect 11886 15722 11942 16000
rect 13450 15722 13506 16000
rect 11886 15694 12388 15722
rect 11886 15600 11942 15694
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4436 14612 4488 14618
rect 4436 14554 4488 14560
rect 4632 14482 4660 14758
rect 5644 14618 5672 15600
rect 5951 15260 6259 15269
rect 5951 15258 5957 15260
rect 6013 15258 6037 15260
rect 6093 15258 6117 15260
rect 6173 15258 6197 15260
rect 6253 15258 6259 15260
rect 6013 15206 6015 15258
rect 6195 15206 6197 15258
rect 5951 15204 5957 15206
rect 6013 15204 6037 15206
rect 6093 15204 6117 15206
rect 6173 15204 6197 15206
rect 6253 15204 6259 15206
rect 5951 15195 6259 15204
rect 7208 14618 7236 15600
rect 8772 15162 8800 15600
rect 9653 15260 9961 15269
rect 9653 15258 9659 15260
rect 9715 15258 9739 15260
rect 9795 15258 9819 15260
rect 9875 15258 9899 15260
rect 9955 15258 9961 15260
rect 9715 15206 9717 15258
rect 9897 15206 9899 15258
rect 9653 15204 9659 15206
rect 9715 15204 9739 15206
rect 9795 15204 9819 15206
rect 9875 15204 9899 15206
rect 9955 15204 9961 15206
rect 9653 15195 9961 15204
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 7802 14716 8110 14725
rect 7802 14714 7808 14716
rect 7864 14714 7888 14716
rect 7944 14714 7968 14716
rect 8024 14714 8048 14716
rect 8104 14714 8110 14716
rect 7864 14662 7866 14714
rect 8046 14662 8048 14714
rect 7802 14660 7808 14662
rect 7864 14660 7888 14662
rect 7944 14660 7968 14662
rect 8024 14660 8048 14662
rect 8104 14660 8110 14662
rect 7802 14651 8110 14660
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 7196 14612 7248 14618
rect 7196 14554 7248 14560
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 5816 14476 5868 14482
rect 5816 14418 5868 14424
rect 6276 14476 6328 14482
rect 6276 14418 6328 14424
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 4100 13628 4408 13637
rect 4100 13626 4106 13628
rect 4162 13626 4186 13628
rect 4242 13626 4266 13628
rect 4322 13626 4346 13628
rect 4402 13626 4408 13628
rect 4162 13574 4164 13626
rect 4344 13574 4346 13626
rect 4100 13572 4106 13574
rect 4162 13572 4186 13574
rect 4242 13572 4266 13574
rect 4322 13572 4346 13574
rect 4402 13572 4408 13574
rect 4100 13563 4408 13572
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3056 13320 3108 13326
rect 3056 13262 3108 13268
rect 2686 12336 2742 12345
rect 2686 12271 2742 12280
rect 3068 12238 3096 13262
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12374 3832 13126
rect 4100 12540 4408 12549
rect 4100 12538 4106 12540
rect 4162 12538 4186 12540
rect 4242 12538 4266 12540
rect 4322 12538 4346 12540
rect 4402 12538 4408 12540
rect 4162 12486 4164 12538
rect 4344 12486 4346 12538
rect 4100 12484 4106 12486
rect 4162 12484 4186 12486
rect 4242 12484 4266 12486
rect 4322 12484 4346 12486
rect 4402 12484 4408 12486
rect 4100 12475 4408 12484
rect 3792 12368 3844 12374
rect 3792 12310 3844 12316
rect 4436 12368 4488 12374
rect 4436 12310 4488 12316
rect 3056 12232 3108 12238
rect 3056 12174 3108 12180
rect 2249 11996 2557 12005
rect 2249 11994 2255 11996
rect 2311 11994 2335 11996
rect 2391 11994 2415 11996
rect 2471 11994 2495 11996
rect 2551 11994 2557 11996
rect 2311 11942 2313 11994
rect 2493 11942 2495 11994
rect 2249 11940 2255 11942
rect 2311 11940 2335 11942
rect 2391 11940 2415 11942
rect 2471 11940 2495 11942
rect 2551 11940 2557 11942
rect 2249 11931 2557 11940
rect 4100 11452 4408 11461
rect 4100 11450 4106 11452
rect 4162 11450 4186 11452
rect 4242 11450 4266 11452
rect 4322 11450 4346 11452
rect 4402 11450 4408 11452
rect 4162 11398 4164 11450
rect 4344 11398 4346 11450
rect 4100 11396 4106 11398
rect 4162 11396 4186 11398
rect 4242 11396 4266 11398
rect 4322 11396 4346 11398
rect 4402 11396 4408 11398
rect 4100 11387 4408 11396
rect 4448 11286 4476 12310
rect 4632 11694 4660 14418
rect 4896 14408 4948 14414
rect 4896 14350 4948 14356
rect 4908 13938 4936 14350
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 4804 13184 4856 13190
rect 4804 13126 4856 13132
rect 4816 12850 4844 13126
rect 4908 12986 4936 13874
rect 5644 13802 5672 14214
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 5184 13326 5212 13398
rect 5552 13394 5580 13670
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 4988 13320 5040 13326
rect 4988 13262 5040 13268
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5000 12986 5028 13262
rect 5184 13190 5212 13262
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 4804 12844 4856 12850
rect 4804 12786 4856 12792
rect 4908 12442 4936 12922
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4724 11898 4752 12310
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 5552 11694 5580 13330
rect 5828 13326 5856 14418
rect 5951 14172 6259 14181
rect 5951 14170 5957 14172
rect 6013 14170 6037 14172
rect 6093 14170 6117 14172
rect 6173 14170 6197 14172
rect 6253 14170 6259 14172
rect 6013 14118 6015 14170
rect 6195 14118 6197 14170
rect 5951 14116 5957 14118
rect 6013 14116 6037 14118
rect 6093 14116 6117 14118
rect 6173 14116 6197 14118
rect 6253 14116 6259 14118
rect 5951 14107 6259 14116
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6196 13530 6224 13738
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5632 12844 5684 12850
rect 5632 12786 5684 12792
rect 5644 11694 5672 12786
rect 5736 12374 5764 13262
rect 5828 12442 5856 13262
rect 5951 13084 6259 13093
rect 5951 13082 5957 13084
rect 6013 13082 6037 13084
rect 6093 13082 6117 13084
rect 6173 13082 6197 13084
rect 6253 13082 6259 13084
rect 6013 13030 6015 13082
rect 6195 13030 6197 13082
rect 5951 13028 5957 13030
rect 6013 13028 6037 13030
rect 6093 13028 6117 13030
rect 6173 13028 6197 13030
rect 6253 13028 6259 13030
rect 5951 13019 6259 13028
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6104 12646 6132 12922
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 5816 12436 5868 12442
rect 5816 12378 5868 12384
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 6104 12306 6132 12582
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 6092 12300 6144 12306
rect 6092 12242 6144 12248
rect 5828 11830 5856 12242
rect 5951 11996 6259 12005
rect 5951 11994 5957 11996
rect 6013 11994 6037 11996
rect 6093 11994 6117 11996
rect 6173 11994 6197 11996
rect 6253 11994 6259 11996
rect 6013 11942 6015 11994
rect 6195 11942 6197 11994
rect 5951 11940 5957 11942
rect 6013 11940 6037 11942
rect 6093 11940 6117 11942
rect 6173 11940 6197 11942
rect 6253 11940 6259 11942
rect 5951 11931 6259 11940
rect 5816 11824 5868 11830
rect 5816 11766 5868 11772
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5632 11688 5684 11694
rect 5632 11630 5684 11636
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 4160 11280 4212 11286
rect 4160 11222 4212 11228
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 2249 10908 2557 10917
rect 2249 10906 2255 10908
rect 2311 10906 2335 10908
rect 2391 10906 2415 10908
rect 2471 10906 2495 10908
rect 2551 10906 2557 10908
rect 2311 10854 2313 10906
rect 2493 10854 2495 10906
rect 2249 10852 2255 10854
rect 2311 10852 2335 10854
rect 2391 10852 2415 10854
rect 2471 10852 2495 10854
rect 2551 10852 2557 10854
rect 2249 10843 2557 10852
rect 4172 10674 4200 11222
rect 5368 11150 5396 11494
rect 6288 11354 6316 14418
rect 6380 14074 6408 14418
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6552 14000 6604 14006
rect 6552 13942 6604 13948
rect 6564 13410 6592 13942
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6472 13382 6592 13410
rect 6932 13410 6960 13670
rect 7024 13530 7052 14350
rect 7116 14074 7144 14486
rect 7760 14074 7788 14486
rect 8208 14340 8260 14346
rect 8208 14282 8260 14288
rect 7104 14068 7156 14074
rect 7104 14010 7156 14016
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7116 13546 7144 14010
rect 8220 14006 8248 14282
rect 8496 14278 8524 14894
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 8484 14272 8536 14278
rect 8484 14214 8536 14220
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8496 13938 8524 14214
rect 8484 13932 8536 13938
rect 8484 13874 8536 13880
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7012 13524 7064 13530
rect 7116 13518 7328 13546
rect 7012 13466 7064 13472
rect 6932 13394 7236 13410
rect 6736 13388 6788 13394
rect 6472 13258 6500 13382
rect 6736 13330 6788 13336
rect 6932 13388 7248 13394
rect 6932 13382 7196 13388
rect 6460 13252 6512 13258
rect 6460 13194 6512 13200
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6472 12481 6500 12650
rect 6458 12472 6514 12481
rect 6458 12407 6514 12416
rect 6564 12374 6592 13194
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6656 12306 6684 13126
rect 6748 12442 6776 13330
rect 6932 13190 6960 13382
rect 7196 13330 7248 13336
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7024 12986 7052 13262
rect 7012 12980 7064 12986
rect 7012 12922 7064 12928
rect 6736 12436 6788 12442
rect 6736 12378 6788 12384
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6380 11830 6408 12106
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 6380 11694 6408 11766
rect 6564 11694 6592 12174
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6276 11348 6328 11354
rect 6276 11290 6328 11296
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5951 10908 6259 10917
rect 5951 10906 5957 10908
rect 6013 10906 6037 10908
rect 6093 10906 6117 10908
rect 6173 10906 6197 10908
rect 6253 10906 6259 10908
rect 6013 10854 6015 10906
rect 6195 10854 6197 10906
rect 5951 10852 5957 10854
rect 6013 10852 6037 10854
rect 6093 10852 6117 10854
rect 6173 10852 6197 10854
rect 6253 10852 6259 10854
rect 5951 10843 6259 10852
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 4100 10364 4408 10373
rect 4100 10362 4106 10364
rect 4162 10362 4186 10364
rect 4242 10362 4266 10364
rect 4322 10362 4346 10364
rect 4402 10362 4408 10364
rect 4162 10310 4164 10362
rect 4344 10310 4346 10362
rect 4100 10308 4106 10310
rect 4162 10308 4186 10310
rect 4242 10308 4266 10310
rect 4322 10308 4346 10310
rect 4402 10308 4408 10310
rect 4100 10299 4408 10308
rect 6288 10266 6316 10542
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 2249 9820 2557 9829
rect 2249 9818 2255 9820
rect 2311 9818 2335 9820
rect 2391 9818 2415 9820
rect 2471 9818 2495 9820
rect 2551 9818 2557 9820
rect 2311 9766 2313 9818
rect 2493 9766 2495 9818
rect 2249 9764 2255 9766
rect 2311 9764 2335 9766
rect 2391 9764 2415 9766
rect 2471 9764 2495 9766
rect 2551 9764 2557 9766
rect 2249 9755 2557 9764
rect 5951 9820 6259 9829
rect 5951 9818 5957 9820
rect 6013 9818 6037 9820
rect 6093 9818 6117 9820
rect 6173 9818 6197 9820
rect 6253 9818 6259 9820
rect 6013 9766 6015 9818
rect 6195 9766 6197 9818
rect 5951 9764 5957 9766
rect 6013 9764 6037 9766
rect 6093 9764 6117 9766
rect 6173 9764 6197 9766
rect 6253 9764 6259 9766
rect 5951 9755 6259 9764
rect 6656 9518 6684 11630
rect 6840 11354 6868 11630
rect 6932 11558 6960 12242
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7300 11218 7328 13518
rect 7668 13394 7696 13670
rect 7802 13628 8110 13637
rect 7802 13626 7808 13628
rect 7864 13626 7888 13628
rect 7944 13626 7968 13628
rect 8024 13626 8048 13628
rect 8104 13626 8110 13628
rect 7864 13574 7866 13626
rect 8046 13574 8048 13626
rect 7802 13572 7808 13574
rect 7864 13572 7888 13574
rect 7944 13572 7968 13574
rect 8024 13572 8048 13574
rect 8104 13572 8110 13574
rect 7802 13563 8110 13572
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7564 13320 7616 13326
rect 7564 13262 7616 13268
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7484 12918 7512 13194
rect 7472 12912 7524 12918
rect 7472 12854 7524 12860
rect 7576 12238 7604 13262
rect 8220 13190 8248 13806
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8392 13320 8444 13326
rect 8392 13262 8444 13268
rect 7656 13184 7708 13190
rect 7656 13126 7708 13132
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 7668 12442 7696 13126
rect 8404 12782 8432 13262
rect 8496 12918 8524 13670
rect 9048 13530 9076 14350
rect 9653 14172 9961 14181
rect 9653 14170 9659 14172
rect 9715 14170 9739 14172
rect 9795 14170 9819 14172
rect 9875 14170 9899 14172
rect 9955 14170 9961 14172
rect 9715 14118 9717 14170
rect 9897 14118 9899 14170
rect 9653 14116 9659 14118
rect 9715 14116 9739 14118
rect 9795 14116 9819 14118
rect 9875 14116 9899 14118
rect 9955 14116 9961 14118
rect 9653 14107 9961 14116
rect 10336 14074 10364 15600
rect 11504 14716 11812 14725
rect 11504 14714 11510 14716
rect 11566 14714 11590 14716
rect 11646 14714 11670 14716
rect 11726 14714 11750 14716
rect 11806 14714 11812 14716
rect 11566 14662 11568 14714
rect 11748 14662 11750 14714
rect 11504 14660 11510 14662
rect 11566 14660 11590 14662
rect 11646 14660 11670 14662
rect 11726 14660 11750 14662
rect 11806 14660 11812 14662
rect 11504 14651 11812 14660
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10968 14476 11020 14482
rect 10968 14418 11020 14424
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9864 13796 9916 13802
rect 9864 13738 9916 13744
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 9128 13388 9180 13394
rect 9232 13376 9260 13738
rect 9180 13348 9260 13376
rect 9128 13330 9180 13336
rect 8484 12912 8536 12918
rect 8484 12854 8536 12860
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8208 12708 8260 12714
rect 8208 12650 8260 12656
rect 7802 12540 8110 12549
rect 7802 12538 7808 12540
rect 7864 12538 7888 12540
rect 7944 12538 7968 12540
rect 8024 12538 8048 12540
rect 8104 12538 8110 12540
rect 7864 12486 7866 12538
rect 8046 12486 8048 12538
rect 7802 12484 7808 12486
rect 7864 12484 7888 12486
rect 7944 12484 7968 12486
rect 8024 12484 8048 12486
rect 8104 12484 8110 12486
rect 7802 12475 8110 12484
rect 8220 12458 8248 12650
rect 7656 12436 7708 12442
rect 8220 12430 8340 12458
rect 7656 12378 7708 12384
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7576 11898 7604 12174
rect 8220 12102 8248 12242
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8312 11898 8340 12430
rect 8404 12102 8432 12718
rect 8496 12442 8524 12854
rect 8588 12782 8616 13330
rect 9232 13190 9260 13348
rect 9312 13320 9364 13326
rect 9312 13262 9364 13268
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 8760 12980 8812 12986
rect 8760 12922 8812 12928
rect 8576 12776 8628 12782
rect 8576 12718 8628 12724
rect 8772 12442 8800 12922
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 6932 10538 6960 11018
rect 7024 10606 7052 11154
rect 7392 11150 7420 11494
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6932 9654 6960 9998
rect 7392 9926 7420 11086
rect 7668 10674 7696 11630
rect 7802 11452 8110 11461
rect 7802 11450 7808 11452
rect 7864 11450 7888 11452
rect 7944 11450 7968 11452
rect 8024 11450 8048 11452
rect 8104 11450 8110 11452
rect 7864 11398 7866 11450
rect 8046 11398 8048 11450
rect 7802 11396 7808 11398
rect 7864 11396 7888 11398
rect 7944 11396 7968 11398
rect 8024 11396 8048 11398
rect 8104 11396 8110 11398
rect 7802 11387 8110 11396
rect 8496 11150 8524 12378
rect 8576 12368 8628 12374
rect 8576 12310 8628 12316
rect 8588 11218 8616 12310
rect 8956 12306 8984 12718
rect 8944 12300 8996 12306
rect 8944 12242 8996 12248
rect 9232 12186 9260 13126
rect 9324 12374 9352 13262
rect 9876 13258 9904 13738
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10152 13394 10180 13466
rect 9956 13388 10008 13394
rect 9956 13330 10008 13336
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 10140 13388 10192 13394
rect 10140 13330 10192 13336
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9968 13190 9996 13330
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9653 13084 9961 13093
rect 9653 13082 9659 13084
rect 9715 13082 9739 13084
rect 9795 13082 9819 13084
rect 9875 13082 9899 13084
rect 9955 13082 9961 13084
rect 9715 13030 9717 13082
rect 9897 13030 9899 13082
rect 9653 13028 9659 13030
rect 9715 13028 9739 13030
rect 9795 13028 9819 13030
rect 9875 13028 9899 13030
rect 9955 13028 9961 13030
rect 9653 13019 9961 13028
rect 10060 12866 10088 13330
rect 9876 12838 10088 12866
rect 9876 12782 9904 12838
rect 9680 12776 9732 12782
rect 9680 12718 9732 12724
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9312 12368 9364 12374
rect 9312 12310 9364 12316
rect 9692 12306 9720 12718
rect 10152 12714 10180 13330
rect 10336 13326 10364 14010
rect 10520 13870 10548 14214
rect 10692 14000 10744 14006
rect 10692 13942 10744 13948
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10704 13394 10732 13942
rect 10796 13870 10824 14418
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10704 13190 10732 13330
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 10048 12232 10100 12238
rect 9232 12158 9352 12186
rect 10048 12174 10100 12180
rect 9324 12102 9352 12158
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 7656 10668 7708 10674
rect 7656 10610 7708 10616
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 7802 10364 8110 10373
rect 7802 10362 7808 10364
rect 7864 10362 7888 10364
rect 7944 10362 7968 10364
rect 8024 10362 8048 10364
rect 8104 10362 8110 10364
rect 7864 10310 7866 10362
rect 8046 10310 8048 10362
rect 7802 10308 7808 10310
rect 7864 10308 7888 10310
rect 7944 10308 7968 10310
rect 8024 10308 8048 10310
rect 8104 10308 8110 10310
rect 7802 10299 8110 10308
rect 8220 10198 8248 10406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 7380 9920 7432 9926
rect 7380 9862 7432 9868
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 7392 9518 7420 9862
rect 8404 9586 8432 10406
rect 8392 9580 8444 9586
rect 8392 9522 8444 9528
rect 6644 9512 6696 9518
rect 6644 9454 6696 9460
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 4100 9276 4408 9285
rect 4100 9274 4106 9276
rect 4162 9274 4186 9276
rect 4242 9274 4266 9276
rect 4322 9274 4346 9276
rect 4402 9274 4408 9276
rect 4162 9222 4164 9274
rect 4344 9222 4346 9274
rect 4100 9220 4106 9222
rect 4162 9220 4186 9222
rect 4242 9220 4266 9222
rect 4322 9220 4346 9222
rect 4402 9220 4408 9222
rect 4100 9211 4408 9220
rect 7802 9276 8110 9285
rect 7802 9274 7808 9276
rect 7864 9274 7888 9276
rect 7944 9274 7968 9276
rect 8024 9274 8048 9276
rect 8104 9274 8110 9276
rect 7864 9222 7866 9274
rect 8046 9222 8048 9274
rect 7802 9220 7808 9222
rect 7864 9220 7888 9222
rect 7944 9220 7968 9222
rect 8024 9220 8048 9222
rect 8104 9220 8110 9222
rect 7802 9211 8110 9220
rect 2249 8732 2557 8741
rect 2249 8730 2255 8732
rect 2311 8730 2335 8732
rect 2391 8730 2415 8732
rect 2471 8730 2495 8732
rect 2551 8730 2557 8732
rect 2311 8678 2313 8730
rect 2493 8678 2495 8730
rect 2249 8676 2255 8678
rect 2311 8676 2335 8678
rect 2391 8676 2415 8678
rect 2471 8676 2495 8678
rect 2551 8676 2557 8678
rect 2249 8667 2557 8676
rect 5951 8732 6259 8741
rect 5951 8730 5957 8732
rect 6013 8730 6037 8732
rect 6093 8730 6117 8732
rect 6173 8730 6197 8732
rect 6253 8730 6259 8732
rect 6013 8678 6015 8730
rect 6195 8678 6197 8730
rect 5951 8676 5957 8678
rect 6013 8676 6037 8678
rect 6093 8676 6117 8678
rect 6173 8676 6197 8678
rect 6253 8676 6259 8678
rect 5951 8667 6259 8676
rect 4100 8188 4408 8197
rect 4100 8186 4106 8188
rect 4162 8186 4186 8188
rect 4242 8186 4266 8188
rect 4322 8186 4346 8188
rect 4402 8186 4408 8188
rect 4162 8134 4164 8186
rect 4344 8134 4346 8186
rect 4100 8132 4106 8134
rect 4162 8132 4186 8134
rect 4242 8132 4266 8134
rect 4322 8132 4346 8134
rect 4402 8132 4408 8134
rect 4100 8123 4408 8132
rect 7802 8188 8110 8197
rect 7802 8186 7808 8188
rect 7864 8186 7888 8188
rect 7944 8186 7968 8188
rect 8024 8186 8048 8188
rect 8104 8186 8110 8188
rect 7864 8134 7866 8186
rect 8046 8134 8048 8186
rect 7802 8132 7808 8134
rect 7864 8132 7888 8134
rect 7944 8132 7968 8134
rect 8024 8132 8048 8134
rect 8104 8132 8110 8134
rect 7802 8123 8110 8132
rect 2249 7644 2557 7653
rect 2249 7642 2255 7644
rect 2311 7642 2335 7644
rect 2391 7642 2415 7644
rect 2471 7642 2495 7644
rect 2551 7642 2557 7644
rect 2311 7590 2313 7642
rect 2493 7590 2495 7642
rect 2249 7588 2255 7590
rect 2311 7588 2335 7590
rect 2391 7588 2415 7590
rect 2471 7588 2495 7590
rect 2551 7588 2557 7590
rect 2249 7579 2557 7588
rect 5951 7644 6259 7653
rect 5951 7642 5957 7644
rect 6013 7642 6037 7644
rect 6093 7642 6117 7644
rect 6173 7642 6197 7644
rect 6253 7642 6259 7644
rect 6013 7590 6015 7642
rect 6195 7590 6197 7642
rect 5951 7588 5957 7590
rect 6013 7588 6037 7590
rect 6093 7588 6117 7590
rect 6173 7588 6197 7590
rect 6253 7588 6259 7590
rect 5951 7579 6259 7588
rect 4100 7100 4408 7109
rect 4100 7098 4106 7100
rect 4162 7098 4186 7100
rect 4242 7098 4266 7100
rect 4322 7098 4346 7100
rect 4402 7098 4408 7100
rect 4162 7046 4164 7098
rect 4344 7046 4346 7098
rect 4100 7044 4106 7046
rect 4162 7044 4186 7046
rect 4242 7044 4266 7046
rect 4322 7044 4346 7046
rect 4402 7044 4408 7046
rect 4100 7035 4408 7044
rect 7802 7100 8110 7109
rect 7802 7098 7808 7100
rect 7864 7098 7888 7100
rect 7944 7098 7968 7100
rect 8024 7098 8048 7100
rect 8104 7098 8110 7100
rect 7864 7046 7866 7098
rect 8046 7046 8048 7098
rect 7802 7044 7808 7046
rect 7864 7044 7888 7046
rect 7944 7044 7968 7046
rect 8024 7044 8048 7046
rect 8104 7044 8110 7046
rect 7802 7035 8110 7044
rect 2249 6556 2557 6565
rect 2249 6554 2255 6556
rect 2311 6554 2335 6556
rect 2391 6554 2415 6556
rect 2471 6554 2495 6556
rect 2551 6554 2557 6556
rect 2311 6502 2313 6554
rect 2493 6502 2495 6554
rect 2249 6500 2255 6502
rect 2311 6500 2335 6502
rect 2391 6500 2415 6502
rect 2471 6500 2495 6502
rect 2551 6500 2557 6502
rect 2249 6491 2557 6500
rect 5951 6556 6259 6565
rect 5951 6554 5957 6556
rect 6013 6554 6037 6556
rect 6093 6554 6117 6556
rect 6173 6554 6197 6556
rect 6253 6554 6259 6556
rect 6013 6502 6015 6554
rect 6195 6502 6197 6554
rect 5951 6500 5957 6502
rect 6013 6500 6037 6502
rect 6093 6500 6117 6502
rect 6173 6500 6197 6502
rect 6253 6500 6259 6502
rect 5951 6491 6259 6500
rect 4100 6012 4408 6021
rect 4100 6010 4106 6012
rect 4162 6010 4186 6012
rect 4242 6010 4266 6012
rect 4322 6010 4346 6012
rect 4402 6010 4408 6012
rect 4162 5958 4164 6010
rect 4344 5958 4346 6010
rect 4100 5956 4106 5958
rect 4162 5956 4186 5958
rect 4242 5956 4266 5958
rect 4322 5956 4346 5958
rect 4402 5956 4408 5958
rect 4100 5947 4408 5956
rect 7802 6012 8110 6021
rect 7802 6010 7808 6012
rect 7864 6010 7888 6012
rect 7944 6010 7968 6012
rect 8024 6010 8048 6012
rect 8104 6010 8110 6012
rect 7864 5958 7866 6010
rect 8046 5958 8048 6010
rect 7802 5956 7808 5958
rect 7864 5956 7888 5958
rect 7944 5956 7968 5958
rect 8024 5956 8048 5958
rect 8104 5956 8110 5958
rect 7802 5947 8110 5956
rect 2249 5468 2557 5477
rect 2249 5466 2255 5468
rect 2311 5466 2335 5468
rect 2391 5466 2415 5468
rect 2471 5466 2495 5468
rect 2551 5466 2557 5468
rect 2311 5414 2313 5466
rect 2493 5414 2495 5466
rect 2249 5412 2255 5414
rect 2311 5412 2335 5414
rect 2391 5412 2415 5414
rect 2471 5412 2495 5414
rect 2551 5412 2557 5414
rect 2249 5403 2557 5412
rect 5951 5468 6259 5477
rect 5951 5466 5957 5468
rect 6013 5466 6037 5468
rect 6093 5466 6117 5468
rect 6173 5466 6197 5468
rect 6253 5466 6259 5468
rect 6013 5414 6015 5466
rect 6195 5414 6197 5466
rect 5951 5412 5957 5414
rect 6013 5412 6037 5414
rect 6093 5412 6117 5414
rect 6173 5412 6197 5414
rect 6253 5412 6259 5414
rect 5951 5403 6259 5412
rect 4100 4924 4408 4933
rect 4100 4922 4106 4924
rect 4162 4922 4186 4924
rect 4242 4922 4266 4924
rect 4322 4922 4346 4924
rect 4402 4922 4408 4924
rect 4162 4870 4164 4922
rect 4344 4870 4346 4922
rect 4100 4868 4106 4870
rect 4162 4868 4186 4870
rect 4242 4868 4266 4870
rect 4322 4868 4346 4870
rect 4402 4868 4408 4870
rect 4100 4859 4408 4868
rect 7802 4924 8110 4933
rect 7802 4922 7808 4924
rect 7864 4922 7888 4924
rect 7944 4922 7968 4924
rect 8024 4922 8048 4924
rect 8104 4922 8110 4924
rect 7864 4870 7866 4922
rect 8046 4870 8048 4922
rect 7802 4868 7808 4870
rect 7864 4868 7888 4870
rect 7944 4868 7968 4870
rect 8024 4868 8048 4870
rect 8104 4868 8110 4870
rect 7802 4859 8110 4868
rect 2249 4380 2557 4389
rect 2249 4378 2255 4380
rect 2311 4378 2335 4380
rect 2391 4378 2415 4380
rect 2471 4378 2495 4380
rect 2551 4378 2557 4380
rect 2311 4326 2313 4378
rect 2493 4326 2495 4378
rect 2249 4324 2255 4326
rect 2311 4324 2335 4326
rect 2391 4324 2415 4326
rect 2471 4324 2495 4326
rect 2551 4324 2557 4326
rect 2249 4315 2557 4324
rect 5951 4380 6259 4389
rect 5951 4378 5957 4380
rect 6013 4378 6037 4380
rect 6093 4378 6117 4380
rect 6173 4378 6197 4380
rect 6253 4378 6259 4380
rect 6013 4326 6015 4378
rect 6195 4326 6197 4378
rect 5951 4324 5957 4326
rect 6013 4324 6037 4326
rect 6093 4324 6117 4326
rect 6173 4324 6197 4326
rect 6253 4324 6259 4326
rect 5951 4315 6259 4324
rect 4100 3836 4408 3845
rect 4100 3834 4106 3836
rect 4162 3834 4186 3836
rect 4242 3834 4266 3836
rect 4322 3834 4346 3836
rect 4402 3834 4408 3836
rect 4162 3782 4164 3834
rect 4344 3782 4346 3834
rect 4100 3780 4106 3782
rect 4162 3780 4186 3782
rect 4242 3780 4266 3782
rect 4322 3780 4346 3782
rect 4402 3780 4408 3782
rect 4100 3771 4408 3780
rect 7802 3836 8110 3845
rect 7802 3834 7808 3836
rect 7864 3834 7888 3836
rect 7944 3834 7968 3836
rect 8024 3834 8048 3836
rect 8104 3834 8110 3836
rect 7864 3782 7866 3834
rect 8046 3782 8048 3834
rect 7802 3780 7808 3782
rect 7864 3780 7888 3782
rect 7944 3780 7968 3782
rect 8024 3780 8048 3782
rect 8104 3780 8110 3782
rect 7802 3771 8110 3780
rect 2249 3292 2557 3301
rect 2249 3290 2255 3292
rect 2311 3290 2335 3292
rect 2391 3290 2415 3292
rect 2471 3290 2495 3292
rect 2551 3290 2557 3292
rect 2311 3238 2313 3290
rect 2493 3238 2495 3290
rect 2249 3236 2255 3238
rect 2311 3236 2335 3238
rect 2391 3236 2415 3238
rect 2471 3236 2495 3238
rect 2551 3236 2557 3238
rect 2249 3227 2557 3236
rect 5951 3292 6259 3301
rect 5951 3290 5957 3292
rect 6013 3290 6037 3292
rect 6093 3290 6117 3292
rect 6173 3290 6197 3292
rect 6253 3290 6259 3292
rect 6013 3238 6015 3290
rect 6195 3238 6197 3290
rect 5951 3236 5957 3238
rect 6013 3236 6037 3238
rect 6093 3236 6117 3238
rect 6173 3236 6197 3238
rect 6253 3236 6259 3238
rect 5951 3227 6259 3236
rect 8680 2774 8708 11222
rect 9048 11218 9076 11290
rect 9140 11218 9168 11494
rect 9324 11286 9352 12038
rect 9653 11996 9961 12005
rect 9653 11994 9659 11996
rect 9715 11994 9739 11996
rect 9795 11994 9819 11996
rect 9875 11994 9899 11996
rect 9955 11994 9961 11996
rect 9715 11942 9717 11994
rect 9897 11942 9899 11994
rect 9653 11940 9659 11942
rect 9715 11940 9739 11942
rect 9795 11940 9819 11942
rect 9875 11940 9899 11942
rect 9955 11940 9961 11942
rect 9653 11931 9961 11940
rect 10060 11898 10088 12174
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9956 11620 10008 11626
rect 9956 11562 10008 11568
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9128 11212 9180 11218
rect 9128 11154 9180 11160
rect 9416 11014 9444 11562
rect 9864 11280 9916 11286
rect 9864 11222 9916 11228
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 8760 11008 8812 11014
rect 8760 10950 8812 10956
rect 9220 11008 9272 11014
rect 9220 10950 9272 10956
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 8772 10130 8800 10950
rect 9232 10606 9260 10950
rect 9508 10810 9536 11154
rect 9876 11014 9904 11222
rect 9968 11218 9996 11562
rect 10152 11234 10180 12650
rect 10244 11830 10272 13126
rect 10796 12986 10824 13330
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 10428 12374 10456 12922
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10152 11218 10272 11234
rect 9956 11212 10008 11218
rect 10152 11212 10284 11218
rect 10152 11206 10232 11212
rect 9956 11154 10008 11160
rect 10232 11154 10284 11160
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 9864 11008 9916 11014
rect 9864 10950 9916 10956
rect 9653 10908 9961 10917
rect 9653 10906 9659 10908
rect 9715 10906 9739 10908
rect 9795 10906 9819 10908
rect 9875 10906 9899 10908
rect 9955 10906 9961 10908
rect 9715 10854 9717 10906
rect 9897 10854 9899 10906
rect 9653 10852 9659 10854
rect 9715 10852 9739 10854
rect 9795 10852 9819 10854
rect 9875 10852 9899 10854
rect 9955 10852 9961 10854
rect 9653 10843 9961 10852
rect 10060 10810 10088 11086
rect 10336 10810 10364 12242
rect 10520 12170 10548 12242
rect 10980 12238 11008 14418
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11256 13530 11284 14350
rect 11808 14074 11836 14486
rect 12360 14278 12388 15694
rect 13096 15694 13506 15722
rect 12348 14272 12400 14278
rect 12348 14214 12400 14220
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 12360 13938 12388 14214
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11348 13394 11376 13670
rect 11504 13628 11812 13637
rect 11504 13626 11510 13628
rect 11566 13626 11590 13628
rect 11646 13626 11670 13628
rect 11726 13626 11750 13628
rect 11806 13626 11812 13628
rect 11566 13574 11568 13626
rect 11748 13574 11750 13626
rect 11504 13572 11510 13574
rect 11566 13572 11590 13574
rect 11646 13572 11670 13574
rect 11726 13572 11750 13574
rect 11806 13572 11812 13574
rect 11504 13563 11812 13572
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 13096 12986 13124 15694
rect 13450 15600 13506 15694
rect 15014 15600 15070 16000
rect 13355 15260 13663 15269
rect 13355 15258 13361 15260
rect 13417 15258 13441 15260
rect 13497 15258 13521 15260
rect 13577 15258 13601 15260
rect 13657 15258 13663 15260
rect 13417 15206 13419 15258
rect 13599 15206 13601 15258
rect 13355 15204 13361 15206
rect 13417 15204 13441 15206
rect 13497 15204 13521 15206
rect 13577 15204 13601 15206
rect 13657 15204 13663 15206
rect 13355 15195 13663 15204
rect 13355 14172 13663 14181
rect 13355 14170 13361 14172
rect 13417 14170 13441 14172
rect 13497 14170 13521 14172
rect 13577 14170 13601 14172
rect 13657 14170 13663 14172
rect 13417 14118 13419 14170
rect 13599 14118 13601 14170
rect 13355 14116 13361 14118
rect 13417 14116 13441 14118
rect 13497 14116 13521 14118
rect 13577 14116 13601 14118
rect 13657 14116 13663 14118
rect 13355 14107 13663 14116
rect 13355 13084 13663 13093
rect 13355 13082 13361 13084
rect 13417 13082 13441 13084
rect 13497 13082 13521 13084
rect 13577 13082 13601 13084
rect 13657 13082 13663 13084
rect 13417 13030 13419 13082
rect 13599 13030 13601 13082
rect 13355 13028 13361 13030
rect 13417 13028 13441 13030
rect 13497 13028 13521 13030
rect 13577 13028 13601 13030
rect 13657 13028 13663 13030
rect 13355 13019 13663 13028
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12716 12776 12768 12782
rect 12716 12718 12768 12724
rect 11504 12540 11812 12549
rect 11504 12538 11510 12540
rect 11566 12538 11590 12540
rect 11646 12538 11670 12540
rect 11726 12538 11750 12540
rect 11806 12538 11812 12540
rect 11566 12486 11568 12538
rect 11748 12486 11750 12538
rect 11504 12484 11510 12486
rect 11566 12484 11590 12486
rect 11646 12484 11670 12486
rect 11726 12484 11750 12486
rect 11806 12484 11812 12486
rect 11504 12475 11812 12484
rect 12728 12442 12756 12718
rect 12716 12436 12768 12442
rect 12716 12378 12768 12384
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10508 12164 10560 12170
rect 10508 12106 10560 12112
rect 10520 11558 10548 12106
rect 10980 11558 11008 12174
rect 12636 11898 12664 12242
rect 12624 11892 12676 11898
rect 12624 11834 12676 11840
rect 13096 11762 13124 12922
rect 13355 11996 13663 12005
rect 13355 11994 13361 11996
rect 13417 11994 13441 11996
rect 13497 11994 13521 11996
rect 13577 11994 13601 11996
rect 13657 11994 13663 11996
rect 13417 11942 13419 11994
rect 13599 11942 13601 11994
rect 13355 11940 13361 11942
rect 13417 11940 13441 11942
rect 13497 11940 13521 11942
rect 13577 11940 13601 11942
rect 13657 11940 13663 11942
rect 13355 11931 13663 11940
rect 15028 11898 15056 15600
rect 15206 14716 15514 14725
rect 15206 14714 15212 14716
rect 15268 14714 15292 14716
rect 15348 14714 15372 14716
rect 15428 14714 15452 14716
rect 15508 14714 15514 14716
rect 15268 14662 15270 14714
rect 15450 14662 15452 14714
rect 15206 14660 15212 14662
rect 15268 14660 15292 14662
rect 15348 14660 15372 14662
rect 15428 14660 15452 14662
rect 15508 14660 15514 14662
rect 15206 14651 15514 14660
rect 15206 13628 15514 13637
rect 15206 13626 15212 13628
rect 15268 13626 15292 13628
rect 15348 13626 15372 13628
rect 15428 13626 15452 13628
rect 15508 13626 15514 13628
rect 15268 13574 15270 13626
rect 15450 13574 15452 13626
rect 15206 13572 15212 13574
rect 15268 13572 15292 13574
rect 15348 13572 15372 13574
rect 15428 13572 15452 13574
rect 15508 13572 15514 13574
rect 15206 13563 15514 13572
rect 15206 12540 15514 12549
rect 15206 12538 15212 12540
rect 15268 12538 15292 12540
rect 15348 12538 15372 12540
rect 15428 12538 15452 12540
rect 15508 12538 15514 12540
rect 15268 12486 15270 12538
rect 15450 12486 15452 12538
rect 15206 12484 15212 12486
rect 15268 12484 15292 12486
rect 15348 12484 15372 12486
rect 15428 12484 15452 12486
rect 15508 12484 15514 12486
rect 15206 12475 15514 12484
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 10508 11552 10560 11558
rect 10508 11494 10560 11500
rect 10968 11552 11020 11558
rect 10968 11494 11020 11500
rect 10520 11218 10548 11494
rect 10508 11212 10560 11218
rect 10508 11154 10560 11160
rect 10980 11150 11008 11494
rect 11504 11452 11812 11461
rect 11504 11450 11510 11452
rect 11566 11450 11590 11452
rect 11646 11450 11670 11452
rect 11726 11450 11750 11452
rect 11806 11450 11812 11452
rect 11566 11398 11568 11450
rect 11748 11398 11750 11450
rect 11504 11396 11510 11398
rect 11566 11396 11590 11398
rect 11646 11396 11670 11398
rect 11726 11396 11750 11398
rect 11806 11396 11812 11398
rect 11504 11387 11812 11396
rect 12176 11354 12204 11630
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10980 10674 11008 11086
rect 11532 10810 11560 11222
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 12544 10606 12572 11630
rect 12728 11354 12756 11630
rect 15206 11452 15514 11461
rect 15206 11450 15212 11452
rect 15268 11450 15292 11452
rect 15348 11450 15372 11452
rect 15428 11450 15452 11452
rect 15508 11450 15514 11452
rect 15268 11398 15270 11450
rect 15450 11398 15452 11450
rect 15206 11396 15212 11398
rect 15268 11396 15292 11398
rect 15348 11396 15372 11398
rect 15428 11396 15452 11398
rect 15508 11396 15514 11398
rect 15206 11387 15514 11396
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 13355 10908 13663 10917
rect 13355 10906 13361 10908
rect 13417 10906 13441 10908
rect 13497 10906 13521 10908
rect 13577 10906 13601 10908
rect 13657 10906 13663 10908
rect 13417 10854 13419 10906
rect 13599 10854 13601 10906
rect 13355 10852 13361 10854
rect 13417 10852 13441 10854
rect 13497 10852 13521 10854
rect 13577 10852 13601 10854
rect 13657 10852 13663 10854
rect 13355 10843 13663 10852
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 9140 10130 9168 10542
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10244 10266 10272 10474
rect 10336 10470 10364 10542
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10336 10130 10364 10406
rect 11504 10364 11812 10373
rect 11504 10362 11510 10364
rect 11566 10362 11590 10364
rect 11646 10362 11670 10364
rect 11726 10362 11750 10364
rect 11806 10362 11812 10364
rect 11566 10310 11568 10362
rect 11748 10310 11750 10362
rect 11504 10308 11510 10310
rect 11566 10308 11590 10310
rect 11646 10308 11670 10310
rect 11726 10308 11750 10310
rect 11806 10308 11812 10310
rect 11504 10299 11812 10308
rect 15206 10364 15514 10373
rect 15206 10362 15212 10364
rect 15268 10362 15292 10364
rect 15348 10362 15372 10364
rect 15428 10362 15452 10364
rect 15508 10362 15514 10364
rect 15268 10310 15270 10362
rect 15450 10310 15452 10362
rect 15206 10308 15212 10310
rect 15268 10308 15292 10310
rect 15348 10308 15372 10310
rect 15428 10308 15452 10310
rect 15508 10308 15514 10310
rect 15206 10299 15514 10308
rect 8760 10124 8812 10130
rect 8760 10066 8812 10072
rect 9128 10124 9180 10130
rect 9128 10066 9180 10072
rect 10324 10124 10376 10130
rect 10324 10066 10376 10072
rect 9653 9820 9961 9829
rect 9653 9818 9659 9820
rect 9715 9818 9739 9820
rect 9795 9818 9819 9820
rect 9875 9818 9899 9820
rect 9955 9818 9961 9820
rect 9715 9766 9717 9818
rect 9897 9766 9899 9818
rect 9653 9764 9659 9766
rect 9715 9764 9739 9766
rect 9795 9764 9819 9766
rect 9875 9764 9899 9766
rect 9955 9764 9961 9766
rect 9653 9755 9961 9764
rect 13355 9820 13663 9829
rect 13355 9818 13361 9820
rect 13417 9818 13441 9820
rect 13497 9818 13521 9820
rect 13577 9818 13601 9820
rect 13657 9818 13663 9820
rect 13417 9766 13419 9818
rect 13599 9766 13601 9818
rect 13355 9764 13361 9766
rect 13417 9764 13441 9766
rect 13497 9764 13521 9766
rect 13577 9764 13601 9766
rect 13657 9764 13663 9766
rect 13355 9755 13663 9764
rect 11504 9276 11812 9285
rect 11504 9274 11510 9276
rect 11566 9274 11590 9276
rect 11646 9274 11670 9276
rect 11726 9274 11750 9276
rect 11806 9274 11812 9276
rect 11566 9222 11568 9274
rect 11748 9222 11750 9274
rect 11504 9220 11510 9222
rect 11566 9220 11590 9222
rect 11646 9220 11670 9222
rect 11726 9220 11750 9222
rect 11806 9220 11812 9222
rect 11504 9211 11812 9220
rect 15206 9276 15514 9285
rect 15206 9274 15212 9276
rect 15268 9274 15292 9276
rect 15348 9274 15372 9276
rect 15428 9274 15452 9276
rect 15508 9274 15514 9276
rect 15268 9222 15270 9274
rect 15450 9222 15452 9274
rect 15206 9220 15212 9222
rect 15268 9220 15292 9222
rect 15348 9220 15372 9222
rect 15428 9220 15452 9222
rect 15508 9220 15514 9222
rect 15206 9211 15514 9220
rect 9653 8732 9961 8741
rect 9653 8730 9659 8732
rect 9715 8730 9739 8732
rect 9795 8730 9819 8732
rect 9875 8730 9899 8732
rect 9955 8730 9961 8732
rect 9715 8678 9717 8730
rect 9897 8678 9899 8730
rect 9653 8676 9659 8678
rect 9715 8676 9739 8678
rect 9795 8676 9819 8678
rect 9875 8676 9899 8678
rect 9955 8676 9961 8678
rect 9653 8667 9961 8676
rect 13355 8732 13663 8741
rect 13355 8730 13361 8732
rect 13417 8730 13441 8732
rect 13497 8730 13521 8732
rect 13577 8730 13601 8732
rect 13657 8730 13663 8732
rect 13417 8678 13419 8730
rect 13599 8678 13601 8730
rect 13355 8676 13361 8678
rect 13417 8676 13441 8678
rect 13497 8676 13521 8678
rect 13577 8676 13601 8678
rect 13657 8676 13663 8678
rect 13355 8667 13663 8676
rect 11504 8188 11812 8197
rect 11504 8186 11510 8188
rect 11566 8186 11590 8188
rect 11646 8186 11670 8188
rect 11726 8186 11750 8188
rect 11806 8186 11812 8188
rect 11566 8134 11568 8186
rect 11748 8134 11750 8186
rect 11504 8132 11510 8134
rect 11566 8132 11590 8134
rect 11646 8132 11670 8134
rect 11726 8132 11750 8134
rect 11806 8132 11812 8134
rect 11504 8123 11812 8132
rect 15206 8188 15514 8197
rect 15206 8186 15212 8188
rect 15268 8186 15292 8188
rect 15348 8186 15372 8188
rect 15428 8186 15452 8188
rect 15508 8186 15514 8188
rect 15268 8134 15270 8186
rect 15450 8134 15452 8186
rect 15206 8132 15212 8134
rect 15268 8132 15292 8134
rect 15348 8132 15372 8134
rect 15428 8132 15452 8134
rect 15508 8132 15514 8134
rect 15206 8123 15514 8132
rect 9653 7644 9961 7653
rect 9653 7642 9659 7644
rect 9715 7642 9739 7644
rect 9795 7642 9819 7644
rect 9875 7642 9899 7644
rect 9955 7642 9961 7644
rect 9715 7590 9717 7642
rect 9897 7590 9899 7642
rect 9653 7588 9659 7590
rect 9715 7588 9739 7590
rect 9795 7588 9819 7590
rect 9875 7588 9899 7590
rect 9955 7588 9961 7590
rect 9653 7579 9961 7588
rect 13355 7644 13663 7653
rect 13355 7642 13361 7644
rect 13417 7642 13441 7644
rect 13497 7642 13521 7644
rect 13577 7642 13601 7644
rect 13657 7642 13663 7644
rect 13417 7590 13419 7642
rect 13599 7590 13601 7642
rect 13355 7588 13361 7590
rect 13417 7588 13441 7590
rect 13497 7588 13521 7590
rect 13577 7588 13601 7590
rect 13657 7588 13663 7590
rect 13355 7579 13663 7588
rect 11504 7100 11812 7109
rect 11504 7098 11510 7100
rect 11566 7098 11590 7100
rect 11646 7098 11670 7100
rect 11726 7098 11750 7100
rect 11806 7098 11812 7100
rect 11566 7046 11568 7098
rect 11748 7046 11750 7098
rect 11504 7044 11510 7046
rect 11566 7044 11590 7046
rect 11646 7044 11670 7046
rect 11726 7044 11750 7046
rect 11806 7044 11812 7046
rect 11504 7035 11812 7044
rect 15206 7100 15514 7109
rect 15206 7098 15212 7100
rect 15268 7098 15292 7100
rect 15348 7098 15372 7100
rect 15428 7098 15452 7100
rect 15508 7098 15514 7100
rect 15268 7046 15270 7098
rect 15450 7046 15452 7098
rect 15206 7044 15212 7046
rect 15268 7044 15292 7046
rect 15348 7044 15372 7046
rect 15428 7044 15452 7046
rect 15508 7044 15514 7046
rect 15206 7035 15514 7044
rect 9653 6556 9961 6565
rect 9653 6554 9659 6556
rect 9715 6554 9739 6556
rect 9795 6554 9819 6556
rect 9875 6554 9899 6556
rect 9955 6554 9961 6556
rect 9715 6502 9717 6554
rect 9897 6502 9899 6554
rect 9653 6500 9659 6502
rect 9715 6500 9739 6502
rect 9795 6500 9819 6502
rect 9875 6500 9899 6502
rect 9955 6500 9961 6502
rect 9653 6491 9961 6500
rect 13355 6556 13663 6565
rect 13355 6554 13361 6556
rect 13417 6554 13441 6556
rect 13497 6554 13521 6556
rect 13577 6554 13601 6556
rect 13657 6554 13663 6556
rect 13417 6502 13419 6554
rect 13599 6502 13601 6554
rect 13355 6500 13361 6502
rect 13417 6500 13441 6502
rect 13497 6500 13521 6502
rect 13577 6500 13601 6502
rect 13657 6500 13663 6502
rect 13355 6491 13663 6500
rect 11504 6012 11812 6021
rect 11504 6010 11510 6012
rect 11566 6010 11590 6012
rect 11646 6010 11670 6012
rect 11726 6010 11750 6012
rect 11806 6010 11812 6012
rect 11566 5958 11568 6010
rect 11748 5958 11750 6010
rect 11504 5956 11510 5958
rect 11566 5956 11590 5958
rect 11646 5956 11670 5958
rect 11726 5956 11750 5958
rect 11806 5956 11812 5958
rect 11504 5947 11812 5956
rect 15206 6012 15514 6021
rect 15206 6010 15212 6012
rect 15268 6010 15292 6012
rect 15348 6010 15372 6012
rect 15428 6010 15452 6012
rect 15508 6010 15514 6012
rect 15268 5958 15270 6010
rect 15450 5958 15452 6010
rect 15206 5956 15212 5958
rect 15268 5956 15292 5958
rect 15348 5956 15372 5958
rect 15428 5956 15452 5958
rect 15508 5956 15514 5958
rect 15206 5947 15514 5956
rect 9653 5468 9961 5477
rect 9653 5466 9659 5468
rect 9715 5466 9739 5468
rect 9795 5466 9819 5468
rect 9875 5466 9899 5468
rect 9955 5466 9961 5468
rect 9715 5414 9717 5466
rect 9897 5414 9899 5466
rect 9653 5412 9659 5414
rect 9715 5412 9739 5414
rect 9795 5412 9819 5414
rect 9875 5412 9899 5414
rect 9955 5412 9961 5414
rect 9653 5403 9961 5412
rect 13355 5468 13663 5477
rect 13355 5466 13361 5468
rect 13417 5466 13441 5468
rect 13497 5466 13521 5468
rect 13577 5466 13601 5468
rect 13657 5466 13663 5468
rect 13417 5414 13419 5466
rect 13599 5414 13601 5466
rect 13355 5412 13361 5414
rect 13417 5412 13441 5414
rect 13497 5412 13521 5414
rect 13577 5412 13601 5414
rect 13657 5412 13663 5414
rect 13355 5403 13663 5412
rect 11504 4924 11812 4933
rect 11504 4922 11510 4924
rect 11566 4922 11590 4924
rect 11646 4922 11670 4924
rect 11726 4922 11750 4924
rect 11806 4922 11812 4924
rect 11566 4870 11568 4922
rect 11748 4870 11750 4922
rect 11504 4868 11510 4870
rect 11566 4868 11590 4870
rect 11646 4868 11670 4870
rect 11726 4868 11750 4870
rect 11806 4868 11812 4870
rect 11504 4859 11812 4868
rect 15206 4924 15514 4933
rect 15206 4922 15212 4924
rect 15268 4922 15292 4924
rect 15348 4922 15372 4924
rect 15428 4922 15452 4924
rect 15508 4922 15514 4924
rect 15268 4870 15270 4922
rect 15450 4870 15452 4922
rect 15206 4868 15212 4870
rect 15268 4868 15292 4870
rect 15348 4868 15372 4870
rect 15428 4868 15452 4870
rect 15508 4868 15514 4870
rect 15206 4859 15514 4868
rect 9653 4380 9961 4389
rect 9653 4378 9659 4380
rect 9715 4378 9739 4380
rect 9795 4378 9819 4380
rect 9875 4378 9899 4380
rect 9955 4378 9961 4380
rect 9715 4326 9717 4378
rect 9897 4326 9899 4378
rect 9653 4324 9659 4326
rect 9715 4324 9739 4326
rect 9795 4324 9819 4326
rect 9875 4324 9899 4326
rect 9955 4324 9961 4326
rect 9653 4315 9961 4324
rect 13355 4380 13663 4389
rect 13355 4378 13361 4380
rect 13417 4378 13441 4380
rect 13497 4378 13521 4380
rect 13577 4378 13601 4380
rect 13657 4378 13663 4380
rect 13417 4326 13419 4378
rect 13599 4326 13601 4378
rect 13355 4324 13361 4326
rect 13417 4324 13441 4326
rect 13497 4324 13521 4326
rect 13577 4324 13601 4326
rect 13657 4324 13663 4326
rect 13355 4315 13663 4324
rect 11504 3836 11812 3845
rect 11504 3834 11510 3836
rect 11566 3834 11590 3836
rect 11646 3834 11670 3836
rect 11726 3834 11750 3836
rect 11806 3834 11812 3836
rect 11566 3782 11568 3834
rect 11748 3782 11750 3834
rect 11504 3780 11510 3782
rect 11566 3780 11590 3782
rect 11646 3780 11670 3782
rect 11726 3780 11750 3782
rect 11806 3780 11812 3782
rect 11504 3771 11812 3780
rect 15206 3836 15514 3845
rect 15206 3834 15212 3836
rect 15268 3834 15292 3836
rect 15348 3834 15372 3836
rect 15428 3834 15452 3836
rect 15508 3834 15514 3836
rect 15268 3782 15270 3834
rect 15450 3782 15452 3834
rect 15206 3780 15212 3782
rect 15268 3780 15292 3782
rect 15348 3780 15372 3782
rect 15428 3780 15452 3782
rect 15508 3780 15514 3782
rect 15206 3771 15514 3780
rect 9653 3292 9961 3301
rect 9653 3290 9659 3292
rect 9715 3290 9739 3292
rect 9795 3290 9819 3292
rect 9875 3290 9899 3292
rect 9955 3290 9961 3292
rect 9715 3238 9717 3290
rect 9897 3238 9899 3290
rect 9653 3236 9659 3238
rect 9715 3236 9739 3238
rect 9795 3236 9819 3238
rect 9875 3236 9899 3238
rect 9955 3236 9961 3238
rect 9653 3227 9961 3236
rect 13355 3292 13663 3301
rect 13355 3290 13361 3292
rect 13417 3290 13441 3292
rect 13497 3290 13521 3292
rect 13577 3290 13601 3292
rect 13657 3290 13663 3292
rect 13417 3238 13419 3290
rect 13599 3238 13601 3290
rect 13355 3236 13361 3238
rect 13417 3236 13441 3238
rect 13497 3236 13521 3238
rect 13577 3236 13601 3238
rect 13657 3236 13663 3238
rect 13355 3227 13663 3236
rect 4100 2748 4408 2757
rect 4100 2746 4106 2748
rect 4162 2746 4186 2748
rect 4242 2746 4266 2748
rect 4322 2746 4346 2748
rect 4402 2746 4408 2748
rect 4162 2694 4164 2746
rect 4344 2694 4346 2746
rect 4100 2692 4106 2694
rect 4162 2692 4186 2694
rect 4242 2692 4266 2694
rect 4322 2692 4346 2694
rect 4402 2692 4408 2694
rect 4100 2683 4408 2692
rect 7802 2748 8110 2757
rect 7802 2746 7808 2748
rect 7864 2746 7888 2748
rect 7944 2746 7968 2748
rect 8024 2746 8048 2748
rect 8104 2746 8110 2748
rect 7864 2694 7866 2746
rect 8046 2694 8048 2746
rect 7802 2692 7808 2694
rect 7864 2692 7888 2694
rect 7944 2692 7968 2694
rect 8024 2692 8048 2694
rect 8104 2692 8110 2694
rect 7802 2683 8110 2692
rect 8588 2746 8708 2774
rect 11504 2748 11812 2757
rect 11504 2746 11510 2748
rect 11566 2746 11590 2748
rect 11646 2746 11670 2748
rect 11726 2746 11750 2748
rect 11806 2746 11812 2748
rect 2249 2204 2557 2213
rect 2249 2202 2255 2204
rect 2311 2202 2335 2204
rect 2391 2202 2415 2204
rect 2471 2202 2495 2204
rect 2551 2202 2557 2204
rect 2311 2150 2313 2202
rect 2493 2150 2495 2202
rect 2249 2148 2255 2150
rect 2311 2148 2335 2150
rect 2391 2148 2415 2150
rect 2471 2148 2495 2150
rect 2551 2148 2557 2150
rect 2249 2139 2557 2148
rect 5951 2204 6259 2213
rect 5951 2202 5957 2204
rect 6013 2202 6037 2204
rect 6093 2202 6117 2204
rect 6173 2202 6197 2204
rect 6253 2202 6259 2204
rect 6013 2150 6015 2202
rect 6195 2150 6197 2202
rect 5951 2148 5957 2150
rect 6013 2148 6037 2150
rect 6093 2148 6117 2150
rect 6173 2148 6197 2150
rect 6253 2148 6259 2150
rect 5951 2139 6259 2148
rect 4100 1660 4408 1669
rect 4100 1658 4106 1660
rect 4162 1658 4186 1660
rect 4242 1658 4266 1660
rect 4322 1658 4346 1660
rect 4402 1658 4408 1660
rect 4162 1606 4164 1658
rect 4344 1606 4346 1658
rect 4100 1604 4106 1606
rect 4162 1604 4186 1606
rect 4242 1604 4266 1606
rect 4322 1604 4346 1606
rect 4402 1604 4408 1606
rect 4100 1595 4408 1604
rect 7802 1660 8110 1669
rect 7802 1658 7808 1660
rect 7864 1658 7888 1660
rect 7944 1658 7968 1660
rect 8024 1658 8048 1660
rect 8104 1658 8110 1660
rect 7864 1606 7866 1658
rect 8046 1606 8048 1658
rect 7802 1604 7808 1606
rect 7864 1604 7888 1606
rect 7944 1604 7968 1606
rect 8024 1604 8048 1606
rect 8104 1604 8110 1606
rect 7802 1595 8110 1604
rect 2249 1116 2557 1125
rect 2249 1114 2255 1116
rect 2311 1114 2335 1116
rect 2391 1114 2415 1116
rect 2471 1114 2495 1116
rect 2551 1114 2557 1116
rect 2311 1062 2313 1114
rect 2493 1062 2495 1114
rect 2249 1060 2255 1062
rect 2311 1060 2335 1062
rect 2391 1060 2415 1062
rect 2471 1060 2495 1062
rect 2551 1060 2557 1062
rect 2249 1051 2557 1060
rect 5951 1116 6259 1125
rect 5951 1114 5957 1116
rect 6013 1114 6037 1116
rect 6093 1114 6117 1116
rect 6173 1114 6197 1116
rect 6253 1114 6259 1116
rect 6013 1062 6015 1114
rect 6195 1062 6197 1114
rect 5951 1060 5957 1062
rect 6013 1060 6037 1062
rect 6093 1060 6117 1062
rect 6173 1060 6197 1062
rect 6253 1060 6259 1062
rect 5951 1051 6259 1060
rect 8588 1018 8616 2746
rect 11566 2694 11568 2746
rect 11748 2694 11750 2746
rect 11504 2692 11510 2694
rect 11566 2692 11590 2694
rect 11646 2692 11670 2694
rect 11726 2692 11750 2694
rect 11806 2692 11812 2694
rect 11504 2683 11812 2692
rect 15206 2748 15514 2757
rect 15206 2746 15212 2748
rect 15268 2746 15292 2748
rect 15348 2746 15372 2748
rect 15428 2746 15452 2748
rect 15508 2746 15514 2748
rect 15268 2694 15270 2746
rect 15450 2694 15452 2746
rect 15206 2692 15212 2694
rect 15268 2692 15292 2694
rect 15348 2692 15372 2694
rect 15428 2692 15452 2694
rect 15508 2692 15514 2694
rect 15206 2683 15514 2692
rect 9653 2204 9961 2213
rect 9653 2202 9659 2204
rect 9715 2202 9739 2204
rect 9795 2202 9819 2204
rect 9875 2202 9899 2204
rect 9955 2202 9961 2204
rect 9715 2150 9717 2202
rect 9897 2150 9899 2202
rect 9653 2148 9659 2150
rect 9715 2148 9739 2150
rect 9795 2148 9819 2150
rect 9875 2148 9899 2150
rect 9955 2148 9961 2150
rect 9653 2139 9961 2148
rect 13355 2204 13663 2213
rect 13355 2202 13361 2204
rect 13417 2202 13441 2204
rect 13497 2202 13521 2204
rect 13577 2202 13601 2204
rect 13657 2202 13663 2204
rect 13417 2150 13419 2202
rect 13599 2150 13601 2202
rect 13355 2148 13361 2150
rect 13417 2148 13441 2150
rect 13497 2148 13521 2150
rect 13577 2148 13601 2150
rect 13657 2148 13663 2150
rect 13355 2139 13663 2148
rect 11504 1660 11812 1669
rect 11504 1658 11510 1660
rect 11566 1658 11590 1660
rect 11646 1658 11670 1660
rect 11726 1658 11750 1660
rect 11806 1658 11812 1660
rect 11566 1606 11568 1658
rect 11748 1606 11750 1658
rect 11504 1604 11510 1606
rect 11566 1604 11590 1606
rect 11646 1604 11670 1606
rect 11726 1604 11750 1606
rect 11806 1604 11812 1606
rect 11504 1595 11812 1604
rect 15206 1660 15514 1669
rect 15206 1658 15212 1660
rect 15268 1658 15292 1660
rect 15348 1658 15372 1660
rect 15428 1658 15452 1660
rect 15508 1658 15514 1660
rect 15268 1606 15270 1658
rect 15450 1606 15452 1658
rect 15206 1604 15212 1606
rect 15268 1604 15292 1606
rect 15348 1604 15372 1606
rect 15428 1604 15452 1606
rect 15508 1604 15514 1606
rect 15206 1595 15514 1604
rect 9653 1116 9961 1125
rect 9653 1114 9659 1116
rect 9715 1114 9739 1116
rect 9795 1114 9819 1116
rect 9875 1114 9899 1116
rect 9955 1114 9961 1116
rect 9715 1062 9717 1114
rect 9897 1062 9899 1114
rect 9653 1060 9659 1062
rect 9715 1060 9739 1062
rect 9795 1060 9819 1062
rect 9875 1060 9899 1062
rect 9955 1060 9961 1062
rect 9653 1051 9961 1060
rect 13355 1116 13663 1125
rect 13355 1114 13361 1116
rect 13417 1114 13441 1116
rect 13497 1114 13521 1116
rect 13577 1114 13601 1116
rect 13657 1114 13663 1116
rect 13417 1062 13419 1114
rect 13599 1062 13601 1114
rect 13355 1060 13361 1062
rect 13417 1060 13441 1062
rect 13497 1060 13521 1062
rect 13577 1060 13601 1062
rect 13657 1060 13663 1062
rect 13355 1051 13663 1060
rect 8576 1012 8628 1018
rect 8576 954 8628 960
rect 8484 740 8536 746
rect 8484 682 8536 688
rect 4100 572 4408 581
rect 4100 570 4106 572
rect 4162 570 4186 572
rect 4242 570 4266 572
rect 4322 570 4346 572
rect 4402 570 4408 572
rect 4162 518 4164 570
rect 4344 518 4346 570
rect 4100 516 4106 518
rect 4162 516 4186 518
rect 4242 516 4266 518
rect 4322 516 4346 518
rect 4402 516 4408 518
rect 4100 507 4408 516
rect 7802 572 8110 581
rect 7802 570 7808 572
rect 7864 570 7888 572
rect 7944 570 7968 572
rect 8024 570 8048 572
rect 8104 570 8110 572
rect 7864 518 7866 570
rect 8046 518 8048 570
rect 7802 516 7808 518
rect 7864 516 7888 518
rect 7944 516 7968 518
rect 8024 516 8048 518
rect 8104 516 8110 518
rect 7802 507 8110 516
rect 8496 474 8524 682
rect 11504 572 11812 581
rect 11504 570 11510 572
rect 11566 570 11590 572
rect 11646 570 11670 572
rect 11726 570 11750 572
rect 11806 570 11812 572
rect 11566 518 11568 570
rect 11748 518 11750 570
rect 11504 516 11510 518
rect 11566 516 11590 518
rect 11646 516 11670 518
rect 11726 516 11750 518
rect 11806 516 11812 518
rect 11504 507 11812 516
rect 15206 572 15514 581
rect 15206 570 15212 572
rect 15268 570 15292 572
rect 15348 570 15372 572
rect 15428 570 15452 572
rect 15508 570 15514 572
rect 15268 518 15270 570
rect 15450 518 15452 570
rect 15206 516 15212 518
rect 15268 516 15292 518
rect 15348 516 15372 518
rect 15428 516 15452 518
rect 15508 516 15514 518
rect 15206 507 15514 516
rect 8024 468 8076 474
rect 7944 428 8024 456
rect 7944 400 7972 428
rect 8024 410 8076 416
rect 8484 468 8536 474
rect 8484 410 8536 416
rect 7930 0 7986 400
<< via2 >>
rect 2255 15258 2311 15260
rect 2335 15258 2391 15260
rect 2415 15258 2471 15260
rect 2495 15258 2551 15260
rect 2255 15206 2301 15258
rect 2301 15206 2311 15258
rect 2335 15206 2365 15258
rect 2365 15206 2377 15258
rect 2377 15206 2391 15258
rect 2415 15206 2429 15258
rect 2429 15206 2441 15258
rect 2441 15206 2471 15258
rect 2495 15206 2505 15258
rect 2505 15206 2551 15258
rect 2255 15204 2311 15206
rect 2335 15204 2391 15206
rect 2415 15204 2471 15206
rect 2495 15204 2551 15206
rect 2255 14170 2311 14172
rect 2335 14170 2391 14172
rect 2415 14170 2471 14172
rect 2495 14170 2551 14172
rect 2255 14118 2301 14170
rect 2301 14118 2311 14170
rect 2335 14118 2365 14170
rect 2365 14118 2377 14170
rect 2377 14118 2391 14170
rect 2415 14118 2429 14170
rect 2429 14118 2441 14170
rect 2441 14118 2471 14170
rect 2495 14118 2505 14170
rect 2505 14118 2551 14170
rect 2255 14116 2311 14118
rect 2335 14116 2391 14118
rect 2415 14116 2471 14118
rect 2495 14116 2551 14118
rect 2255 13082 2311 13084
rect 2335 13082 2391 13084
rect 2415 13082 2471 13084
rect 2495 13082 2551 13084
rect 2255 13030 2301 13082
rect 2301 13030 2311 13082
rect 2335 13030 2365 13082
rect 2365 13030 2377 13082
rect 2377 13030 2391 13082
rect 2415 13030 2429 13082
rect 2429 13030 2441 13082
rect 2441 13030 2471 13082
rect 2495 13030 2505 13082
rect 2505 13030 2551 13082
rect 2255 13028 2311 13030
rect 2335 13028 2391 13030
rect 2415 13028 2471 13030
rect 2495 13028 2551 13030
rect 4106 14714 4162 14716
rect 4186 14714 4242 14716
rect 4266 14714 4322 14716
rect 4346 14714 4402 14716
rect 4106 14662 4152 14714
rect 4152 14662 4162 14714
rect 4186 14662 4216 14714
rect 4216 14662 4228 14714
rect 4228 14662 4242 14714
rect 4266 14662 4280 14714
rect 4280 14662 4292 14714
rect 4292 14662 4322 14714
rect 4346 14662 4356 14714
rect 4356 14662 4402 14714
rect 4106 14660 4162 14662
rect 4186 14660 4242 14662
rect 4266 14660 4322 14662
rect 4346 14660 4402 14662
rect 5957 15258 6013 15260
rect 6037 15258 6093 15260
rect 6117 15258 6173 15260
rect 6197 15258 6253 15260
rect 5957 15206 6003 15258
rect 6003 15206 6013 15258
rect 6037 15206 6067 15258
rect 6067 15206 6079 15258
rect 6079 15206 6093 15258
rect 6117 15206 6131 15258
rect 6131 15206 6143 15258
rect 6143 15206 6173 15258
rect 6197 15206 6207 15258
rect 6207 15206 6253 15258
rect 5957 15204 6013 15206
rect 6037 15204 6093 15206
rect 6117 15204 6173 15206
rect 6197 15204 6253 15206
rect 9659 15258 9715 15260
rect 9739 15258 9795 15260
rect 9819 15258 9875 15260
rect 9899 15258 9955 15260
rect 9659 15206 9705 15258
rect 9705 15206 9715 15258
rect 9739 15206 9769 15258
rect 9769 15206 9781 15258
rect 9781 15206 9795 15258
rect 9819 15206 9833 15258
rect 9833 15206 9845 15258
rect 9845 15206 9875 15258
rect 9899 15206 9909 15258
rect 9909 15206 9955 15258
rect 9659 15204 9715 15206
rect 9739 15204 9795 15206
rect 9819 15204 9875 15206
rect 9899 15204 9955 15206
rect 7808 14714 7864 14716
rect 7888 14714 7944 14716
rect 7968 14714 8024 14716
rect 8048 14714 8104 14716
rect 7808 14662 7854 14714
rect 7854 14662 7864 14714
rect 7888 14662 7918 14714
rect 7918 14662 7930 14714
rect 7930 14662 7944 14714
rect 7968 14662 7982 14714
rect 7982 14662 7994 14714
rect 7994 14662 8024 14714
rect 8048 14662 8058 14714
rect 8058 14662 8104 14714
rect 7808 14660 7864 14662
rect 7888 14660 7944 14662
rect 7968 14660 8024 14662
rect 8048 14660 8104 14662
rect 4106 13626 4162 13628
rect 4186 13626 4242 13628
rect 4266 13626 4322 13628
rect 4346 13626 4402 13628
rect 4106 13574 4152 13626
rect 4152 13574 4162 13626
rect 4186 13574 4216 13626
rect 4216 13574 4228 13626
rect 4228 13574 4242 13626
rect 4266 13574 4280 13626
rect 4280 13574 4292 13626
rect 4292 13574 4322 13626
rect 4346 13574 4356 13626
rect 4356 13574 4402 13626
rect 4106 13572 4162 13574
rect 4186 13572 4242 13574
rect 4266 13572 4322 13574
rect 4346 13572 4402 13574
rect 2686 12280 2742 12336
rect 4106 12538 4162 12540
rect 4186 12538 4242 12540
rect 4266 12538 4322 12540
rect 4346 12538 4402 12540
rect 4106 12486 4152 12538
rect 4152 12486 4162 12538
rect 4186 12486 4216 12538
rect 4216 12486 4228 12538
rect 4228 12486 4242 12538
rect 4266 12486 4280 12538
rect 4280 12486 4292 12538
rect 4292 12486 4322 12538
rect 4346 12486 4356 12538
rect 4356 12486 4402 12538
rect 4106 12484 4162 12486
rect 4186 12484 4242 12486
rect 4266 12484 4322 12486
rect 4346 12484 4402 12486
rect 2255 11994 2311 11996
rect 2335 11994 2391 11996
rect 2415 11994 2471 11996
rect 2495 11994 2551 11996
rect 2255 11942 2301 11994
rect 2301 11942 2311 11994
rect 2335 11942 2365 11994
rect 2365 11942 2377 11994
rect 2377 11942 2391 11994
rect 2415 11942 2429 11994
rect 2429 11942 2441 11994
rect 2441 11942 2471 11994
rect 2495 11942 2505 11994
rect 2505 11942 2551 11994
rect 2255 11940 2311 11942
rect 2335 11940 2391 11942
rect 2415 11940 2471 11942
rect 2495 11940 2551 11942
rect 4106 11450 4162 11452
rect 4186 11450 4242 11452
rect 4266 11450 4322 11452
rect 4346 11450 4402 11452
rect 4106 11398 4152 11450
rect 4152 11398 4162 11450
rect 4186 11398 4216 11450
rect 4216 11398 4228 11450
rect 4228 11398 4242 11450
rect 4266 11398 4280 11450
rect 4280 11398 4292 11450
rect 4292 11398 4322 11450
rect 4346 11398 4356 11450
rect 4356 11398 4402 11450
rect 4106 11396 4162 11398
rect 4186 11396 4242 11398
rect 4266 11396 4322 11398
rect 4346 11396 4402 11398
rect 5957 14170 6013 14172
rect 6037 14170 6093 14172
rect 6117 14170 6173 14172
rect 6197 14170 6253 14172
rect 5957 14118 6003 14170
rect 6003 14118 6013 14170
rect 6037 14118 6067 14170
rect 6067 14118 6079 14170
rect 6079 14118 6093 14170
rect 6117 14118 6131 14170
rect 6131 14118 6143 14170
rect 6143 14118 6173 14170
rect 6197 14118 6207 14170
rect 6207 14118 6253 14170
rect 5957 14116 6013 14118
rect 6037 14116 6093 14118
rect 6117 14116 6173 14118
rect 6197 14116 6253 14118
rect 5957 13082 6013 13084
rect 6037 13082 6093 13084
rect 6117 13082 6173 13084
rect 6197 13082 6253 13084
rect 5957 13030 6003 13082
rect 6003 13030 6013 13082
rect 6037 13030 6067 13082
rect 6067 13030 6079 13082
rect 6079 13030 6093 13082
rect 6117 13030 6131 13082
rect 6131 13030 6143 13082
rect 6143 13030 6173 13082
rect 6197 13030 6207 13082
rect 6207 13030 6253 13082
rect 5957 13028 6013 13030
rect 6037 13028 6093 13030
rect 6117 13028 6173 13030
rect 6197 13028 6253 13030
rect 5957 11994 6013 11996
rect 6037 11994 6093 11996
rect 6117 11994 6173 11996
rect 6197 11994 6253 11996
rect 5957 11942 6003 11994
rect 6003 11942 6013 11994
rect 6037 11942 6067 11994
rect 6067 11942 6079 11994
rect 6079 11942 6093 11994
rect 6117 11942 6131 11994
rect 6131 11942 6143 11994
rect 6143 11942 6173 11994
rect 6197 11942 6207 11994
rect 6207 11942 6253 11994
rect 5957 11940 6013 11942
rect 6037 11940 6093 11942
rect 6117 11940 6173 11942
rect 6197 11940 6253 11942
rect 2255 10906 2311 10908
rect 2335 10906 2391 10908
rect 2415 10906 2471 10908
rect 2495 10906 2551 10908
rect 2255 10854 2301 10906
rect 2301 10854 2311 10906
rect 2335 10854 2365 10906
rect 2365 10854 2377 10906
rect 2377 10854 2391 10906
rect 2415 10854 2429 10906
rect 2429 10854 2441 10906
rect 2441 10854 2471 10906
rect 2495 10854 2505 10906
rect 2505 10854 2551 10906
rect 2255 10852 2311 10854
rect 2335 10852 2391 10854
rect 2415 10852 2471 10854
rect 2495 10852 2551 10854
rect 6458 12416 6514 12472
rect 5957 10906 6013 10908
rect 6037 10906 6093 10908
rect 6117 10906 6173 10908
rect 6197 10906 6253 10908
rect 5957 10854 6003 10906
rect 6003 10854 6013 10906
rect 6037 10854 6067 10906
rect 6067 10854 6079 10906
rect 6079 10854 6093 10906
rect 6117 10854 6131 10906
rect 6131 10854 6143 10906
rect 6143 10854 6173 10906
rect 6197 10854 6207 10906
rect 6207 10854 6253 10906
rect 5957 10852 6013 10854
rect 6037 10852 6093 10854
rect 6117 10852 6173 10854
rect 6197 10852 6253 10854
rect 4106 10362 4162 10364
rect 4186 10362 4242 10364
rect 4266 10362 4322 10364
rect 4346 10362 4402 10364
rect 4106 10310 4152 10362
rect 4152 10310 4162 10362
rect 4186 10310 4216 10362
rect 4216 10310 4228 10362
rect 4228 10310 4242 10362
rect 4266 10310 4280 10362
rect 4280 10310 4292 10362
rect 4292 10310 4322 10362
rect 4346 10310 4356 10362
rect 4356 10310 4402 10362
rect 4106 10308 4162 10310
rect 4186 10308 4242 10310
rect 4266 10308 4322 10310
rect 4346 10308 4402 10310
rect 2255 9818 2311 9820
rect 2335 9818 2391 9820
rect 2415 9818 2471 9820
rect 2495 9818 2551 9820
rect 2255 9766 2301 9818
rect 2301 9766 2311 9818
rect 2335 9766 2365 9818
rect 2365 9766 2377 9818
rect 2377 9766 2391 9818
rect 2415 9766 2429 9818
rect 2429 9766 2441 9818
rect 2441 9766 2471 9818
rect 2495 9766 2505 9818
rect 2505 9766 2551 9818
rect 2255 9764 2311 9766
rect 2335 9764 2391 9766
rect 2415 9764 2471 9766
rect 2495 9764 2551 9766
rect 5957 9818 6013 9820
rect 6037 9818 6093 9820
rect 6117 9818 6173 9820
rect 6197 9818 6253 9820
rect 5957 9766 6003 9818
rect 6003 9766 6013 9818
rect 6037 9766 6067 9818
rect 6067 9766 6079 9818
rect 6079 9766 6093 9818
rect 6117 9766 6131 9818
rect 6131 9766 6143 9818
rect 6143 9766 6173 9818
rect 6197 9766 6207 9818
rect 6207 9766 6253 9818
rect 5957 9764 6013 9766
rect 6037 9764 6093 9766
rect 6117 9764 6173 9766
rect 6197 9764 6253 9766
rect 7808 13626 7864 13628
rect 7888 13626 7944 13628
rect 7968 13626 8024 13628
rect 8048 13626 8104 13628
rect 7808 13574 7854 13626
rect 7854 13574 7864 13626
rect 7888 13574 7918 13626
rect 7918 13574 7930 13626
rect 7930 13574 7944 13626
rect 7968 13574 7982 13626
rect 7982 13574 7994 13626
rect 7994 13574 8024 13626
rect 8048 13574 8058 13626
rect 8058 13574 8104 13626
rect 7808 13572 7864 13574
rect 7888 13572 7944 13574
rect 7968 13572 8024 13574
rect 8048 13572 8104 13574
rect 9659 14170 9715 14172
rect 9739 14170 9795 14172
rect 9819 14170 9875 14172
rect 9899 14170 9955 14172
rect 9659 14118 9705 14170
rect 9705 14118 9715 14170
rect 9739 14118 9769 14170
rect 9769 14118 9781 14170
rect 9781 14118 9795 14170
rect 9819 14118 9833 14170
rect 9833 14118 9845 14170
rect 9845 14118 9875 14170
rect 9899 14118 9909 14170
rect 9909 14118 9955 14170
rect 9659 14116 9715 14118
rect 9739 14116 9795 14118
rect 9819 14116 9875 14118
rect 9899 14116 9955 14118
rect 11510 14714 11566 14716
rect 11590 14714 11646 14716
rect 11670 14714 11726 14716
rect 11750 14714 11806 14716
rect 11510 14662 11556 14714
rect 11556 14662 11566 14714
rect 11590 14662 11620 14714
rect 11620 14662 11632 14714
rect 11632 14662 11646 14714
rect 11670 14662 11684 14714
rect 11684 14662 11696 14714
rect 11696 14662 11726 14714
rect 11750 14662 11760 14714
rect 11760 14662 11806 14714
rect 11510 14660 11566 14662
rect 11590 14660 11646 14662
rect 11670 14660 11726 14662
rect 11750 14660 11806 14662
rect 7808 12538 7864 12540
rect 7888 12538 7944 12540
rect 7968 12538 8024 12540
rect 8048 12538 8104 12540
rect 7808 12486 7854 12538
rect 7854 12486 7864 12538
rect 7888 12486 7918 12538
rect 7918 12486 7930 12538
rect 7930 12486 7944 12538
rect 7968 12486 7982 12538
rect 7982 12486 7994 12538
rect 7994 12486 8024 12538
rect 8048 12486 8058 12538
rect 8058 12486 8104 12538
rect 7808 12484 7864 12486
rect 7888 12484 7944 12486
rect 7968 12484 8024 12486
rect 8048 12484 8104 12486
rect 7808 11450 7864 11452
rect 7888 11450 7944 11452
rect 7968 11450 8024 11452
rect 8048 11450 8104 11452
rect 7808 11398 7854 11450
rect 7854 11398 7864 11450
rect 7888 11398 7918 11450
rect 7918 11398 7930 11450
rect 7930 11398 7944 11450
rect 7968 11398 7982 11450
rect 7982 11398 7994 11450
rect 7994 11398 8024 11450
rect 8048 11398 8058 11450
rect 8058 11398 8104 11450
rect 7808 11396 7864 11398
rect 7888 11396 7944 11398
rect 7968 11396 8024 11398
rect 8048 11396 8104 11398
rect 9659 13082 9715 13084
rect 9739 13082 9795 13084
rect 9819 13082 9875 13084
rect 9899 13082 9955 13084
rect 9659 13030 9705 13082
rect 9705 13030 9715 13082
rect 9739 13030 9769 13082
rect 9769 13030 9781 13082
rect 9781 13030 9795 13082
rect 9819 13030 9833 13082
rect 9833 13030 9845 13082
rect 9845 13030 9875 13082
rect 9899 13030 9909 13082
rect 9909 13030 9955 13082
rect 9659 13028 9715 13030
rect 9739 13028 9795 13030
rect 9819 13028 9875 13030
rect 9899 13028 9955 13030
rect 7808 10362 7864 10364
rect 7888 10362 7944 10364
rect 7968 10362 8024 10364
rect 8048 10362 8104 10364
rect 7808 10310 7854 10362
rect 7854 10310 7864 10362
rect 7888 10310 7918 10362
rect 7918 10310 7930 10362
rect 7930 10310 7944 10362
rect 7968 10310 7982 10362
rect 7982 10310 7994 10362
rect 7994 10310 8024 10362
rect 8048 10310 8058 10362
rect 8058 10310 8104 10362
rect 7808 10308 7864 10310
rect 7888 10308 7944 10310
rect 7968 10308 8024 10310
rect 8048 10308 8104 10310
rect 4106 9274 4162 9276
rect 4186 9274 4242 9276
rect 4266 9274 4322 9276
rect 4346 9274 4402 9276
rect 4106 9222 4152 9274
rect 4152 9222 4162 9274
rect 4186 9222 4216 9274
rect 4216 9222 4228 9274
rect 4228 9222 4242 9274
rect 4266 9222 4280 9274
rect 4280 9222 4292 9274
rect 4292 9222 4322 9274
rect 4346 9222 4356 9274
rect 4356 9222 4402 9274
rect 4106 9220 4162 9222
rect 4186 9220 4242 9222
rect 4266 9220 4322 9222
rect 4346 9220 4402 9222
rect 7808 9274 7864 9276
rect 7888 9274 7944 9276
rect 7968 9274 8024 9276
rect 8048 9274 8104 9276
rect 7808 9222 7854 9274
rect 7854 9222 7864 9274
rect 7888 9222 7918 9274
rect 7918 9222 7930 9274
rect 7930 9222 7944 9274
rect 7968 9222 7982 9274
rect 7982 9222 7994 9274
rect 7994 9222 8024 9274
rect 8048 9222 8058 9274
rect 8058 9222 8104 9274
rect 7808 9220 7864 9222
rect 7888 9220 7944 9222
rect 7968 9220 8024 9222
rect 8048 9220 8104 9222
rect 2255 8730 2311 8732
rect 2335 8730 2391 8732
rect 2415 8730 2471 8732
rect 2495 8730 2551 8732
rect 2255 8678 2301 8730
rect 2301 8678 2311 8730
rect 2335 8678 2365 8730
rect 2365 8678 2377 8730
rect 2377 8678 2391 8730
rect 2415 8678 2429 8730
rect 2429 8678 2441 8730
rect 2441 8678 2471 8730
rect 2495 8678 2505 8730
rect 2505 8678 2551 8730
rect 2255 8676 2311 8678
rect 2335 8676 2391 8678
rect 2415 8676 2471 8678
rect 2495 8676 2551 8678
rect 5957 8730 6013 8732
rect 6037 8730 6093 8732
rect 6117 8730 6173 8732
rect 6197 8730 6253 8732
rect 5957 8678 6003 8730
rect 6003 8678 6013 8730
rect 6037 8678 6067 8730
rect 6067 8678 6079 8730
rect 6079 8678 6093 8730
rect 6117 8678 6131 8730
rect 6131 8678 6143 8730
rect 6143 8678 6173 8730
rect 6197 8678 6207 8730
rect 6207 8678 6253 8730
rect 5957 8676 6013 8678
rect 6037 8676 6093 8678
rect 6117 8676 6173 8678
rect 6197 8676 6253 8678
rect 4106 8186 4162 8188
rect 4186 8186 4242 8188
rect 4266 8186 4322 8188
rect 4346 8186 4402 8188
rect 4106 8134 4152 8186
rect 4152 8134 4162 8186
rect 4186 8134 4216 8186
rect 4216 8134 4228 8186
rect 4228 8134 4242 8186
rect 4266 8134 4280 8186
rect 4280 8134 4292 8186
rect 4292 8134 4322 8186
rect 4346 8134 4356 8186
rect 4356 8134 4402 8186
rect 4106 8132 4162 8134
rect 4186 8132 4242 8134
rect 4266 8132 4322 8134
rect 4346 8132 4402 8134
rect 7808 8186 7864 8188
rect 7888 8186 7944 8188
rect 7968 8186 8024 8188
rect 8048 8186 8104 8188
rect 7808 8134 7854 8186
rect 7854 8134 7864 8186
rect 7888 8134 7918 8186
rect 7918 8134 7930 8186
rect 7930 8134 7944 8186
rect 7968 8134 7982 8186
rect 7982 8134 7994 8186
rect 7994 8134 8024 8186
rect 8048 8134 8058 8186
rect 8058 8134 8104 8186
rect 7808 8132 7864 8134
rect 7888 8132 7944 8134
rect 7968 8132 8024 8134
rect 8048 8132 8104 8134
rect 2255 7642 2311 7644
rect 2335 7642 2391 7644
rect 2415 7642 2471 7644
rect 2495 7642 2551 7644
rect 2255 7590 2301 7642
rect 2301 7590 2311 7642
rect 2335 7590 2365 7642
rect 2365 7590 2377 7642
rect 2377 7590 2391 7642
rect 2415 7590 2429 7642
rect 2429 7590 2441 7642
rect 2441 7590 2471 7642
rect 2495 7590 2505 7642
rect 2505 7590 2551 7642
rect 2255 7588 2311 7590
rect 2335 7588 2391 7590
rect 2415 7588 2471 7590
rect 2495 7588 2551 7590
rect 5957 7642 6013 7644
rect 6037 7642 6093 7644
rect 6117 7642 6173 7644
rect 6197 7642 6253 7644
rect 5957 7590 6003 7642
rect 6003 7590 6013 7642
rect 6037 7590 6067 7642
rect 6067 7590 6079 7642
rect 6079 7590 6093 7642
rect 6117 7590 6131 7642
rect 6131 7590 6143 7642
rect 6143 7590 6173 7642
rect 6197 7590 6207 7642
rect 6207 7590 6253 7642
rect 5957 7588 6013 7590
rect 6037 7588 6093 7590
rect 6117 7588 6173 7590
rect 6197 7588 6253 7590
rect 4106 7098 4162 7100
rect 4186 7098 4242 7100
rect 4266 7098 4322 7100
rect 4346 7098 4402 7100
rect 4106 7046 4152 7098
rect 4152 7046 4162 7098
rect 4186 7046 4216 7098
rect 4216 7046 4228 7098
rect 4228 7046 4242 7098
rect 4266 7046 4280 7098
rect 4280 7046 4292 7098
rect 4292 7046 4322 7098
rect 4346 7046 4356 7098
rect 4356 7046 4402 7098
rect 4106 7044 4162 7046
rect 4186 7044 4242 7046
rect 4266 7044 4322 7046
rect 4346 7044 4402 7046
rect 7808 7098 7864 7100
rect 7888 7098 7944 7100
rect 7968 7098 8024 7100
rect 8048 7098 8104 7100
rect 7808 7046 7854 7098
rect 7854 7046 7864 7098
rect 7888 7046 7918 7098
rect 7918 7046 7930 7098
rect 7930 7046 7944 7098
rect 7968 7046 7982 7098
rect 7982 7046 7994 7098
rect 7994 7046 8024 7098
rect 8048 7046 8058 7098
rect 8058 7046 8104 7098
rect 7808 7044 7864 7046
rect 7888 7044 7944 7046
rect 7968 7044 8024 7046
rect 8048 7044 8104 7046
rect 2255 6554 2311 6556
rect 2335 6554 2391 6556
rect 2415 6554 2471 6556
rect 2495 6554 2551 6556
rect 2255 6502 2301 6554
rect 2301 6502 2311 6554
rect 2335 6502 2365 6554
rect 2365 6502 2377 6554
rect 2377 6502 2391 6554
rect 2415 6502 2429 6554
rect 2429 6502 2441 6554
rect 2441 6502 2471 6554
rect 2495 6502 2505 6554
rect 2505 6502 2551 6554
rect 2255 6500 2311 6502
rect 2335 6500 2391 6502
rect 2415 6500 2471 6502
rect 2495 6500 2551 6502
rect 5957 6554 6013 6556
rect 6037 6554 6093 6556
rect 6117 6554 6173 6556
rect 6197 6554 6253 6556
rect 5957 6502 6003 6554
rect 6003 6502 6013 6554
rect 6037 6502 6067 6554
rect 6067 6502 6079 6554
rect 6079 6502 6093 6554
rect 6117 6502 6131 6554
rect 6131 6502 6143 6554
rect 6143 6502 6173 6554
rect 6197 6502 6207 6554
rect 6207 6502 6253 6554
rect 5957 6500 6013 6502
rect 6037 6500 6093 6502
rect 6117 6500 6173 6502
rect 6197 6500 6253 6502
rect 4106 6010 4162 6012
rect 4186 6010 4242 6012
rect 4266 6010 4322 6012
rect 4346 6010 4402 6012
rect 4106 5958 4152 6010
rect 4152 5958 4162 6010
rect 4186 5958 4216 6010
rect 4216 5958 4228 6010
rect 4228 5958 4242 6010
rect 4266 5958 4280 6010
rect 4280 5958 4292 6010
rect 4292 5958 4322 6010
rect 4346 5958 4356 6010
rect 4356 5958 4402 6010
rect 4106 5956 4162 5958
rect 4186 5956 4242 5958
rect 4266 5956 4322 5958
rect 4346 5956 4402 5958
rect 7808 6010 7864 6012
rect 7888 6010 7944 6012
rect 7968 6010 8024 6012
rect 8048 6010 8104 6012
rect 7808 5958 7854 6010
rect 7854 5958 7864 6010
rect 7888 5958 7918 6010
rect 7918 5958 7930 6010
rect 7930 5958 7944 6010
rect 7968 5958 7982 6010
rect 7982 5958 7994 6010
rect 7994 5958 8024 6010
rect 8048 5958 8058 6010
rect 8058 5958 8104 6010
rect 7808 5956 7864 5958
rect 7888 5956 7944 5958
rect 7968 5956 8024 5958
rect 8048 5956 8104 5958
rect 2255 5466 2311 5468
rect 2335 5466 2391 5468
rect 2415 5466 2471 5468
rect 2495 5466 2551 5468
rect 2255 5414 2301 5466
rect 2301 5414 2311 5466
rect 2335 5414 2365 5466
rect 2365 5414 2377 5466
rect 2377 5414 2391 5466
rect 2415 5414 2429 5466
rect 2429 5414 2441 5466
rect 2441 5414 2471 5466
rect 2495 5414 2505 5466
rect 2505 5414 2551 5466
rect 2255 5412 2311 5414
rect 2335 5412 2391 5414
rect 2415 5412 2471 5414
rect 2495 5412 2551 5414
rect 5957 5466 6013 5468
rect 6037 5466 6093 5468
rect 6117 5466 6173 5468
rect 6197 5466 6253 5468
rect 5957 5414 6003 5466
rect 6003 5414 6013 5466
rect 6037 5414 6067 5466
rect 6067 5414 6079 5466
rect 6079 5414 6093 5466
rect 6117 5414 6131 5466
rect 6131 5414 6143 5466
rect 6143 5414 6173 5466
rect 6197 5414 6207 5466
rect 6207 5414 6253 5466
rect 5957 5412 6013 5414
rect 6037 5412 6093 5414
rect 6117 5412 6173 5414
rect 6197 5412 6253 5414
rect 4106 4922 4162 4924
rect 4186 4922 4242 4924
rect 4266 4922 4322 4924
rect 4346 4922 4402 4924
rect 4106 4870 4152 4922
rect 4152 4870 4162 4922
rect 4186 4870 4216 4922
rect 4216 4870 4228 4922
rect 4228 4870 4242 4922
rect 4266 4870 4280 4922
rect 4280 4870 4292 4922
rect 4292 4870 4322 4922
rect 4346 4870 4356 4922
rect 4356 4870 4402 4922
rect 4106 4868 4162 4870
rect 4186 4868 4242 4870
rect 4266 4868 4322 4870
rect 4346 4868 4402 4870
rect 7808 4922 7864 4924
rect 7888 4922 7944 4924
rect 7968 4922 8024 4924
rect 8048 4922 8104 4924
rect 7808 4870 7854 4922
rect 7854 4870 7864 4922
rect 7888 4870 7918 4922
rect 7918 4870 7930 4922
rect 7930 4870 7944 4922
rect 7968 4870 7982 4922
rect 7982 4870 7994 4922
rect 7994 4870 8024 4922
rect 8048 4870 8058 4922
rect 8058 4870 8104 4922
rect 7808 4868 7864 4870
rect 7888 4868 7944 4870
rect 7968 4868 8024 4870
rect 8048 4868 8104 4870
rect 2255 4378 2311 4380
rect 2335 4378 2391 4380
rect 2415 4378 2471 4380
rect 2495 4378 2551 4380
rect 2255 4326 2301 4378
rect 2301 4326 2311 4378
rect 2335 4326 2365 4378
rect 2365 4326 2377 4378
rect 2377 4326 2391 4378
rect 2415 4326 2429 4378
rect 2429 4326 2441 4378
rect 2441 4326 2471 4378
rect 2495 4326 2505 4378
rect 2505 4326 2551 4378
rect 2255 4324 2311 4326
rect 2335 4324 2391 4326
rect 2415 4324 2471 4326
rect 2495 4324 2551 4326
rect 5957 4378 6013 4380
rect 6037 4378 6093 4380
rect 6117 4378 6173 4380
rect 6197 4378 6253 4380
rect 5957 4326 6003 4378
rect 6003 4326 6013 4378
rect 6037 4326 6067 4378
rect 6067 4326 6079 4378
rect 6079 4326 6093 4378
rect 6117 4326 6131 4378
rect 6131 4326 6143 4378
rect 6143 4326 6173 4378
rect 6197 4326 6207 4378
rect 6207 4326 6253 4378
rect 5957 4324 6013 4326
rect 6037 4324 6093 4326
rect 6117 4324 6173 4326
rect 6197 4324 6253 4326
rect 4106 3834 4162 3836
rect 4186 3834 4242 3836
rect 4266 3834 4322 3836
rect 4346 3834 4402 3836
rect 4106 3782 4152 3834
rect 4152 3782 4162 3834
rect 4186 3782 4216 3834
rect 4216 3782 4228 3834
rect 4228 3782 4242 3834
rect 4266 3782 4280 3834
rect 4280 3782 4292 3834
rect 4292 3782 4322 3834
rect 4346 3782 4356 3834
rect 4356 3782 4402 3834
rect 4106 3780 4162 3782
rect 4186 3780 4242 3782
rect 4266 3780 4322 3782
rect 4346 3780 4402 3782
rect 7808 3834 7864 3836
rect 7888 3834 7944 3836
rect 7968 3834 8024 3836
rect 8048 3834 8104 3836
rect 7808 3782 7854 3834
rect 7854 3782 7864 3834
rect 7888 3782 7918 3834
rect 7918 3782 7930 3834
rect 7930 3782 7944 3834
rect 7968 3782 7982 3834
rect 7982 3782 7994 3834
rect 7994 3782 8024 3834
rect 8048 3782 8058 3834
rect 8058 3782 8104 3834
rect 7808 3780 7864 3782
rect 7888 3780 7944 3782
rect 7968 3780 8024 3782
rect 8048 3780 8104 3782
rect 2255 3290 2311 3292
rect 2335 3290 2391 3292
rect 2415 3290 2471 3292
rect 2495 3290 2551 3292
rect 2255 3238 2301 3290
rect 2301 3238 2311 3290
rect 2335 3238 2365 3290
rect 2365 3238 2377 3290
rect 2377 3238 2391 3290
rect 2415 3238 2429 3290
rect 2429 3238 2441 3290
rect 2441 3238 2471 3290
rect 2495 3238 2505 3290
rect 2505 3238 2551 3290
rect 2255 3236 2311 3238
rect 2335 3236 2391 3238
rect 2415 3236 2471 3238
rect 2495 3236 2551 3238
rect 5957 3290 6013 3292
rect 6037 3290 6093 3292
rect 6117 3290 6173 3292
rect 6197 3290 6253 3292
rect 5957 3238 6003 3290
rect 6003 3238 6013 3290
rect 6037 3238 6067 3290
rect 6067 3238 6079 3290
rect 6079 3238 6093 3290
rect 6117 3238 6131 3290
rect 6131 3238 6143 3290
rect 6143 3238 6173 3290
rect 6197 3238 6207 3290
rect 6207 3238 6253 3290
rect 5957 3236 6013 3238
rect 6037 3236 6093 3238
rect 6117 3236 6173 3238
rect 6197 3236 6253 3238
rect 9659 11994 9715 11996
rect 9739 11994 9795 11996
rect 9819 11994 9875 11996
rect 9899 11994 9955 11996
rect 9659 11942 9705 11994
rect 9705 11942 9715 11994
rect 9739 11942 9769 11994
rect 9769 11942 9781 11994
rect 9781 11942 9795 11994
rect 9819 11942 9833 11994
rect 9833 11942 9845 11994
rect 9845 11942 9875 11994
rect 9899 11942 9909 11994
rect 9909 11942 9955 11994
rect 9659 11940 9715 11942
rect 9739 11940 9795 11942
rect 9819 11940 9875 11942
rect 9899 11940 9955 11942
rect 9659 10906 9715 10908
rect 9739 10906 9795 10908
rect 9819 10906 9875 10908
rect 9899 10906 9955 10908
rect 9659 10854 9705 10906
rect 9705 10854 9715 10906
rect 9739 10854 9769 10906
rect 9769 10854 9781 10906
rect 9781 10854 9795 10906
rect 9819 10854 9833 10906
rect 9833 10854 9845 10906
rect 9845 10854 9875 10906
rect 9899 10854 9909 10906
rect 9909 10854 9955 10906
rect 9659 10852 9715 10854
rect 9739 10852 9795 10854
rect 9819 10852 9875 10854
rect 9899 10852 9955 10854
rect 11510 13626 11566 13628
rect 11590 13626 11646 13628
rect 11670 13626 11726 13628
rect 11750 13626 11806 13628
rect 11510 13574 11556 13626
rect 11556 13574 11566 13626
rect 11590 13574 11620 13626
rect 11620 13574 11632 13626
rect 11632 13574 11646 13626
rect 11670 13574 11684 13626
rect 11684 13574 11696 13626
rect 11696 13574 11726 13626
rect 11750 13574 11760 13626
rect 11760 13574 11806 13626
rect 11510 13572 11566 13574
rect 11590 13572 11646 13574
rect 11670 13572 11726 13574
rect 11750 13572 11806 13574
rect 13361 15258 13417 15260
rect 13441 15258 13497 15260
rect 13521 15258 13577 15260
rect 13601 15258 13657 15260
rect 13361 15206 13407 15258
rect 13407 15206 13417 15258
rect 13441 15206 13471 15258
rect 13471 15206 13483 15258
rect 13483 15206 13497 15258
rect 13521 15206 13535 15258
rect 13535 15206 13547 15258
rect 13547 15206 13577 15258
rect 13601 15206 13611 15258
rect 13611 15206 13657 15258
rect 13361 15204 13417 15206
rect 13441 15204 13497 15206
rect 13521 15204 13577 15206
rect 13601 15204 13657 15206
rect 13361 14170 13417 14172
rect 13441 14170 13497 14172
rect 13521 14170 13577 14172
rect 13601 14170 13657 14172
rect 13361 14118 13407 14170
rect 13407 14118 13417 14170
rect 13441 14118 13471 14170
rect 13471 14118 13483 14170
rect 13483 14118 13497 14170
rect 13521 14118 13535 14170
rect 13535 14118 13547 14170
rect 13547 14118 13577 14170
rect 13601 14118 13611 14170
rect 13611 14118 13657 14170
rect 13361 14116 13417 14118
rect 13441 14116 13497 14118
rect 13521 14116 13577 14118
rect 13601 14116 13657 14118
rect 13361 13082 13417 13084
rect 13441 13082 13497 13084
rect 13521 13082 13577 13084
rect 13601 13082 13657 13084
rect 13361 13030 13407 13082
rect 13407 13030 13417 13082
rect 13441 13030 13471 13082
rect 13471 13030 13483 13082
rect 13483 13030 13497 13082
rect 13521 13030 13535 13082
rect 13535 13030 13547 13082
rect 13547 13030 13577 13082
rect 13601 13030 13611 13082
rect 13611 13030 13657 13082
rect 13361 13028 13417 13030
rect 13441 13028 13497 13030
rect 13521 13028 13577 13030
rect 13601 13028 13657 13030
rect 11510 12538 11566 12540
rect 11590 12538 11646 12540
rect 11670 12538 11726 12540
rect 11750 12538 11806 12540
rect 11510 12486 11556 12538
rect 11556 12486 11566 12538
rect 11590 12486 11620 12538
rect 11620 12486 11632 12538
rect 11632 12486 11646 12538
rect 11670 12486 11684 12538
rect 11684 12486 11696 12538
rect 11696 12486 11726 12538
rect 11750 12486 11760 12538
rect 11760 12486 11806 12538
rect 11510 12484 11566 12486
rect 11590 12484 11646 12486
rect 11670 12484 11726 12486
rect 11750 12484 11806 12486
rect 13361 11994 13417 11996
rect 13441 11994 13497 11996
rect 13521 11994 13577 11996
rect 13601 11994 13657 11996
rect 13361 11942 13407 11994
rect 13407 11942 13417 11994
rect 13441 11942 13471 11994
rect 13471 11942 13483 11994
rect 13483 11942 13497 11994
rect 13521 11942 13535 11994
rect 13535 11942 13547 11994
rect 13547 11942 13577 11994
rect 13601 11942 13611 11994
rect 13611 11942 13657 11994
rect 13361 11940 13417 11942
rect 13441 11940 13497 11942
rect 13521 11940 13577 11942
rect 13601 11940 13657 11942
rect 15212 14714 15268 14716
rect 15292 14714 15348 14716
rect 15372 14714 15428 14716
rect 15452 14714 15508 14716
rect 15212 14662 15258 14714
rect 15258 14662 15268 14714
rect 15292 14662 15322 14714
rect 15322 14662 15334 14714
rect 15334 14662 15348 14714
rect 15372 14662 15386 14714
rect 15386 14662 15398 14714
rect 15398 14662 15428 14714
rect 15452 14662 15462 14714
rect 15462 14662 15508 14714
rect 15212 14660 15268 14662
rect 15292 14660 15348 14662
rect 15372 14660 15428 14662
rect 15452 14660 15508 14662
rect 15212 13626 15268 13628
rect 15292 13626 15348 13628
rect 15372 13626 15428 13628
rect 15452 13626 15508 13628
rect 15212 13574 15258 13626
rect 15258 13574 15268 13626
rect 15292 13574 15322 13626
rect 15322 13574 15334 13626
rect 15334 13574 15348 13626
rect 15372 13574 15386 13626
rect 15386 13574 15398 13626
rect 15398 13574 15428 13626
rect 15452 13574 15462 13626
rect 15462 13574 15508 13626
rect 15212 13572 15268 13574
rect 15292 13572 15348 13574
rect 15372 13572 15428 13574
rect 15452 13572 15508 13574
rect 15212 12538 15268 12540
rect 15292 12538 15348 12540
rect 15372 12538 15428 12540
rect 15452 12538 15508 12540
rect 15212 12486 15258 12538
rect 15258 12486 15268 12538
rect 15292 12486 15322 12538
rect 15322 12486 15334 12538
rect 15334 12486 15348 12538
rect 15372 12486 15386 12538
rect 15386 12486 15398 12538
rect 15398 12486 15428 12538
rect 15452 12486 15462 12538
rect 15462 12486 15508 12538
rect 15212 12484 15268 12486
rect 15292 12484 15348 12486
rect 15372 12484 15428 12486
rect 15452 12484 15508 12486
rect 11510 11450 11566 11452
rect 11590 11450 11646 11452
rect 11670 11450 11726 11452
rect 11750 11450 11806 11452
rect 11510 11398 11556 11450
rect 11556 11398 11566 11450
rect 11590 11398 11620 11450
rect 11620 11398 11632 11450
rect 11632 11398 11646 11450
rect 11670 11398 11684 11450
rect 11684 11398 11696 11450
rect 11696 11398 11726 11450
rect 11750 11398 11760 11450
rect 11760 11398 11806 11450
rect 11510 11396 11566 11398
rect 11590 11396 11646 11398
rect 11670 11396 11726 11398
rect 11750 11396 11806 11398
rect 15212 11450 15268 11452
rect 15292 11450 15348 11452
rect 15372 11450 15428 11452
rect 15452 11450 15508 11452
rect 15212 11398 15258 11450
rect 15258 11398 15268 11450
rect 15292 11398 15322 11450
rect 15322 11398 15334 11450
rect 15334 11398 15348 11450
rect 15372 11398 15386 11450
rect 15386 11398 15398 11450
rect 15398 11398 15428 11450
rect 15452 11398 15462 11450
rect 15462 11398 15508 11450
rect 15212 11396 15268 11398
rect 15292 11396 15348 11398
rect 15372 11396 15428 11398
rect 15452 11396 15508 11398
rect 13361 10906 13417 10908
rect 13441 10906 13497 10908
rect 13521 10906 13577 10908
rect 13601 10906 13657 10908
rect 13361 10854 13407 10906
rect 13407 10854 13417 10906
rect 13441 10854 13471 10906
rect 13471 10854 13483 10906
rect 13483 10854 13497 10906
rect 13521 10854 13535 10906
rect 13535 10854 13547 10906
rect 13547 10854 13577 10906
rect 13601 10854 13611 10906
rect 13611 10854 13657 10906
rect 13361 10852 13417 10854
rect 13441 10852 13497 10854
rect 13521 10852 13577 10854
rect 13601 10852 13657 10854
rect 11510 10362 11566 10364
rect 11590 10362 11646 10364
rect 11670 10362 11726 10364
rect 11750 10362 11806 10364
rect 11510 10310 11556 10362
rect 11556 10310 11566 10362
rect 11590 10310 11620 10362
rect 11620 10310 11632 10362
rect 11632 10310 11646 10362
rect 11670 10310 11684 10362
rect 11684 10310 11696 10362
rect 11696 10310 11726 10362
rect 11750 10310 11760 10362
rect 11760 10310 11806 10362
rect 11510 10308 11566 10310
rect 11590 10308 11646 10310
rect 11670 10308 11726 10310
rect 11750 10308 11806 10310
rect 15212 10362 15268 10364
rect 15292 10362 15348 10364
rect 15372 10362 15428 10364
rect 15452 10362 15508 10364
rect 15212 10310 15258 10362
rect 15258 10310 15268 10362
rect 15292 10310 15322 10362
rect 15322 10310 15334 10362
rect 15334 10310 15348 10362
rect 15372 10310 15386 10362
rect 15386 10310 15398 10362
rect 15398 10310 15428 10362
rect 15452 10310 15462 10362
rect 15462 10310 15508 10362
rect 15212 10308 15268 10310
rect 15292 10308 15348 10310
rect 15372 10308 15428 10310
rect 15452 10308 15508 10310
rect 9659 9818 9715 9820
rect 9739 9818 9795 9820
rect 9819 9818 9875 9820
rect 9899 9818 9955 9820
rect 9659 9766 9705 9818
rect 9705 9766 9715 9818
rect 9739 9766 9769 9818
rect 9769 9766 9781 9818
rect 9781 9766 9795 9818
rect 9819 9766 9833 9818
rect 9833 9766 9845 9818
rect 9845 9766 9875 9818
rect 9899 9766 9909 9818
rect 9909 9766 9955 9818
rect 9659 9764 9715 9766
rect 9739 9764 9795 9766
rect 9819 9764 9875 9766
rect 9899 9764 9955 9766
rect 13361 9818 13417 9820
rect 13441 9818 13497 9820
rect 13521 9818 13577 9820
rect 13601 9818 13657 9820
rect 13361 9766 13407 9818
rect 13407 9766 13417 9818
rect 13441 9766 13471 9818
rect 13471 9766 13483 9818
rect 13483 9766 13497 9818
rect 13521 9766 13535 9818
rect 13535 9766 13547 9818
rect 13547 9766 13577 9818
rect 13601 9766 13611 9818
rect 13611 9766 13657 9818
rect 13361 9764 13417 9766
rect 13441 9764 13497 9766
rect 13521 9764 13577 9766
rect 13601 9764 13657 9766
rect 11510 9274 11566 9276
rect 11590 9274 11646 9276
rect 11670 9274 11726 9276
rect 11750 9274 11806 9276
rect 11510 9222 11556 9274
rect 11556 9222 11566 9274
rect 11590 9222 11620 9274
rect 11620 9222 11632 9274
rect 11632 9222 11646 9274
rect 11670 9222 11684 9274
rect 11684 9222 11696 9274
rect 11696 9222 11726 9274
rect 11750 9222 11760 9274
rect 11760 9222 11806 9274
rect 11510 9220 11566 9222
rect 11590 9220 11646 9222
rect 11670 9220 11726 9222
rect 11750 9220 11806 9222
rect 15212 9274 15268 9276
rect 15292 9274 15348 9276
rect 15372 9274 15428 9276
rect 15452 9274 15508 9276
rect 15212 9222 15258 9274
rect 15258 9222 15268 9274
rect 15292 9222 15322 9274
rect 15322 9222 15334 9274
rect 15334 9222 15348 9274
rect 15372 9222 15386 9274
rect 15386 9222 15398 9274
rect 15398 9222 15428 9274
rect 15452 9222 15462 9274
rect 15462 9222 15508 9274
rect 15212 9220 15268 9222
rect 15292 9220 15348 9222
rect 15372 9220 15428 9222
rect 15452 9220 15508 9222
rect 9659 8730 9715 8732
rect 9739 8730 9795 8732
rect 9819 8730 9875 8732
rect 9899 8730 9955 8732
rect 9659 8678 9705 8730
rect 9705 8678 9715 8730
rect 9739 8678 9769 8730
rect 9769 8678 9781 8730
rect 9781 8678 9795 8730
rect 9819 8678 9833 8730
rect 9833 8678 9845 8730
rect 9845 8678 9875 8730
rect 9899 8678 9909 8730
rect 9909 8678 9955 8730
rect 9659 8676 9715 8678
rect 9739 8676 9795 8678
rect 9819 8676 9875 8678
rect 9899 8676 9955 8678
rect 13361 8730 13417 8732
rect 13441 8730 13497 8732
rect 13521 8730 13577 8732
rect 13601 8730 13657 8732
rect 13361 8678 13407 8730
rect 13407 8678 13417 8730
rect 13441 8678 13471 8730
rect 13471 8678 13483 8730
rect 13483 8678 13497 8730
rect 13521 8678 13535 8730
rect 13535 8678 13547 8730
rect 13547 8678 13577 8730
rect 13601 8678 13611 8730
rect 13611 8678 13657 8730
rect 13361 8676 13417 8678
rect 13441 8676 13497 8678
rect 13521 8676 13577 8678
rect 13601 8676 13657 8678
rect 11510 8186 11566 8188
rect 11590 8186 11646 8188
rect 11670 8186 11726 8188
rect 11750 8186 11806 8188
rect 11510 8134 11556 8186
rect 11556 8134 11566 8186
rect 11590 8134 11620 8186
rect 11620 8134 11632 8186
rect 11632 8134 11646 8186
rect 11670 8134 11684 8186
rect 11684 8134 11696 8186
rect 11696 8134 11726 8186
rect 11750 8134 11760 8186
rect 11760 8134 11806 8186
rect 11510 8132 11566 8134
rect 11590 8132 11646 8134
rect 11670 8132 11726 8134
rect 11750 8132 11806 8134
rect 15212 8186 15268 8188
rect 15292 8186 15348 8188
rect 15372 8186 15428 8188
rect 15452 8186 15508 8188
rect 15212 8134 15258 8186
rect 15258 8134 15268 8186
rect 15292 8134 15322 8186
rect 15322 8134 15334 8186
rect 15334 8134 15348 8186
rect 15372 8134 15386 8186
rect 15386 8134 15398 8186
rect 15398 8134 15428 8186
rect 15452 8134 15462 8186
rect 15462 8134 15508 8186
rect 15212 8132 15268 8134
rect 15292 8132 15348 8134
rect 15372 8132 15428 8134
rect 15452 8132 15508 8134
rect 9659 7642 9715 7644
rect 9739 7642 9795 7644
rect 9819 7642 9875 7644
rect 9899 7642 9955 7644
rect 9659 7590 9705 7642
rect 9705 7590 9715 7642
rect 9739 7590 9769 7642
rect 9769 7590 9781 7642
rect 9781 7590 9795 7642
rect 9819 7590 9833 7642
rect 9833 7590 9845 7642
rect 9845 7590 9875 7642
rect 9899 7590 9909 7642
rect 9909 7590 9955 7642
rect 9659 7588 9715 7590
rect 9739 7588 9795 7590
rect 9819 7588 9875 7590
rect 9899 7588 9955 7590
rect 13361 7642 13417 7644
rect 13441 7642 13497 7644
rect 13521 7642 13577 7644
rect 13601 7642 13657 7644
rect 13361 7590 13407 7642
rect 13407 7590 13417 7642
rect 13441 7590 13471 7642
rect 13471 7590 13483 7642
rect 13483 7590 13497 7642
rect 13521 7590 13535 7642
rect 13535 7590 13547 7642
rect 13547 7590 13577 7642
rect 13601 7590 13611 7642
rect 13611 7590 13657 7642
rect 13361 7588 13417 7590
rect 13441 7588 13497 7590
rect 13521 7588 13577 7590
rect 13601 7588 13657 7590
rect 11510 7098 11566 7100
rect 11590 7098 11646 7100
rect 11670 7098 11726 7100
rect 11750 7098 11806 7100
rect 11510 7046 11556 7098
rect 11556 7046 11566 7098
rect 11590 7046 11620 7098
rect 11620 7046 11632 7098
rect 11632 7046 11646 7098
rect 11670 7046 11684 7098
rect 11684 7046 11696 7098
rect 11696 7046 11726 7098
rect 11750 7046 11760 7098
rect 11760 7046 11806 7098
rect 11510 7044 11566 7046
rect 11590 7044 11646 7046
rect 11670 7044 11726 7046
rect 11750 7044 11806 7046
rect 15212 7098 15268 7100
rect 15292 7098 15348 7100
rect 15372 7098 15428 7100
rect 15452 7098 15508 7100
rect 15212 7046 15258 7098
rect 15258 7046 15268 7098
rect 15292 7046 15322 7098
rect 15322 7046 15334 7098
rect 15334 7046 15348 7098
rect 15372 7046 15386 7098
rect 15386 7046 15398 7098
rect 15398 7046 15428 7098
rect 15452 7046 15462 7098
rect 15462 7046 15508 7098
rect 15212 7044 15268 7046
rect 15292 7044 15348 7046
rect 15372 7044 15428 7046
rect 15452 7044 15508 7046
rect 9659 6554 9715 6556
rect 9739 6554 9795 6556
rect 9819 6554 9875 6556
rect 9899 6554 9955 6556
rect 9659 6502 9705 6554
rect 9705 6502 9715 6554
rect 9739 6502 9769 6554
rect 9769 6502 9781 6554
rect 9781 6502 9795 6554
rect 9819 6502 9833 6554
rect 9833 6502 9845 6554
rect 9845 6502 9875 6554
rect 9899 6502 9909 6554
rect 9909 6502 9955 6554
rect 9659 6500 9715 6502
rect 9739 6500 9795 6502
rect 9819 6500 9875 6502
rect 9899 6500 9955 6502
rect 13361 6554 13417 6556
rect 13441 6554 13497 6556
rect 13521 6554 13577 6556
rect 13601 6554 13657 6556
rect 13361 6502 13407 6554
rect 13407 6502 13417 6554
rect 13441 6502 13471 6554
rect 13471 6502 13483 6554
rect 13483 6502 13497 6554
rect 13521 6502 13535 6554
rect 13535 6502 13547 6554
rect 13547 6502 13577 6554
rect 13601 6502 13611 6554
rect 13611 6502 13657 6554
rect 13361 6500 13417 6502
rect 13441 6500 13497 6502
rect 13521 6500 13577 6502
rect 13601 6500 13657 6502
rect 11510 6010 11566 6012
rect 11590 6010 11646 6012
rect 11670 6010 11726 6012
rect 11750 6010 11806 6012
rect 11510 5958 11556 6010
rect 11556 5958 11566 6010
rect 11590 5958 11620 6010
rect 11620 5958 11632 6010
rect 11632 5958 11646 6010
rect 11670 5958 11684 6010
rect 11684 5958 11696 6010
rect 11696 5958 11726 6010
rect 11750 5958 11760 6010
rect 11760 5958 11806 6010
rect 11510 5956 11566 5958
rect 11590 5956 11646 5958
rect 11670 5956 11726 5958
rect 11750 5956 11806 5958
rect 15212 6010 15268 6012
rect 15292 6010 15348 6012
rect 15372 6010 15428 6012
rect 15452 6010 15508 6012
rect 15212 5958 15258 6010
rect 15258 5958 15268 6010
rect 15292 5958 15322 6010
rect 15322 5958 15334 6010
rect 15334 5958 15348 6010
rect 15372 5958 15386 6010
rect 15386 5958 15398 6010
rect 15398 5958 15428 6010
rect 15452 5958 15462 6010
rect 15462 5958 15508 6010
rect 15212 5956 15268 5958
rect 15292 5956 15348 5958
rect 15372 5956 15428 5958
rect 15452 5956 15508 5958
rect 9659 5466 9715 5468
rect 9739 5466 9795 5468
rect 9819 5466 9875 5468
rect 9899 5466 9955 5468
rect 9659 5414 9705 5466
rect 9705 5414 9715 5466
rect 9739 5414 9769 5466
rect 9769 5414 9781 5466
rect 9781 5414 9795 5466
rect 9819 5414 9833 5466
rect 9833 5414 9845 5466
rect 9845 5414 9875 5466
rect 9899 5414 9909 5466
rect 9909 5414 9955 5466
rect 9659 5412 9715 5414
rect 9739 5412 9795 5414
rect 9819 5412 9875 5414
rect 9899 5412 9955 5414
rect 13361 5466 13417 5468
rect 13441 5466 13497 5468
rect 13521 5466 13577 5468
rect 13601 5466 13657 5468
rect 13361 5414 13407 5466
rect 13407 5414 13417 5466
rect 13441 5414 13471 5466
rect 13471 5414 13483 5466
rect 13483 5414 13497 5466
rect 13521 5414 13535 5466
rect 13535 5414 13547 5466
rect 13547 5414 13577 5466
rect 13601 5414 13611 5466
rect 13611 5414 13657 5466
rect 13361 5412 13417 5414
rect 13441 5412 13497 5414
rect 13521 5412 13577 5414
rect 13601 5412 13657 5414
rect 11510 4922 11566 4924
rect 11590 4922 11646 4924
rect 11670 4922 11726 4924
rect 11750 4922 11806 4924
rect 11510 4870 11556 4922
rect 11556 4870 11566 4922
rect 11590 4870 11620 4922
rect 11620 4870 11632 4922
rect 11632 4870 11646 4922
rect 11670 4870 11684 4922
rect 11684 4870 11696 4922
rect 11696 4870 11726 4922
rect 11750 4870 11760 4922
rect 11760 4870 11806 4922
rect 11510 4868 11566 4870
rect 11590 4868 11646 4870
rect 11670 4868 11726 4870
rect 11750 4868 11806 4870
rect 15212 4922 15268 4924
rect 15292 4922 15348 4924
rect 15372 4922 15428 4924
rect 15452 4922 15508 4924
rect 15212 4870 15258 4922
rect 15258 4870 15268 4922
rect 15292 4870 15322 4922
rect 15322 4870 15334 4922
rect 15334 4870 15348 4922
rect 15372 4870 15386 4922
rect 15386 4870 15398 4922
rect 15398 4870 15428 4922
rect 15452 4870 15462 4922
rect 15462 4870 15508 4922
rect 15212 4868 15268 4870
rect 15292 4868 15348 4870
rect 15372 4868 15428 4870
rect 15452 4868 15508 4870
rect 9659 4378 9715 4380
rect 9739 4378 9795 4380
rect 9819 4378 9875 4380
rect 9899 4378 9955 4380
rect 9659 4326 9705 4378
rect 9705 4326 9715 4378
rect 9739 4326 9769 4378
rect 9769 4326 9781 4378
rect 9781 4326 9795 4378
rect 9819 4326 9833 4378
rect 9833 4326 9845 4378
rect 9845 4326 9875 4378
rect 9899 4326 9909 4378
rect 9909 4326 9955 4378
rect 9659 4324 9715 4326
rect 9739 4324 9795 4326
rect 9819 4324 9875 4326
rect 9899 4324 9955 4326
rect 13361 4378 13417 4380
rect 13441 4378 13497 4380
rect 13521 4378 13577 4380
rect 13601 4378 13657 4380
rect 13361 4326 13407 4378
rect 13407 4326 13417 4378
rect 13441 4326 13471 4378
rect 13471 4326 13483 4378
rect 13483 4326 13497 4378
rect 13521 4326 13535 4378
rect 13535 4326 13547 4378
rect 13547 4326 13577 4378
rect 13601 4326 13611 4378
rect 13611 4326 13657 4378
rect 13361 4324 13417 4326
rect 13441 4324 13497 4326
rect 13521 4324 13577 4326
rect 13601 4324 13657 4326
rect 11510 3834 11566 3836
rect 11590 3834 11646 3836
rect 11670 3834 11726 3836
rect 11750 3834 11806 3836
rect 11510 3782 11556 3834
rect 11556 3782 11566 3834
rect 11590 3782 11620 3834
rect 11620 3782 11632 3834
rect 11632 3782 11646 3834
rect 11670 3782 11684 3834
rect 11684 3782 11696 3834
rect 11696 3782 11726 3834
rect 11750 3782 11760 3834
rect 11760 3782 11806 3834
rect 11510 3780 11566 3782
rect 11590 3780 11646 3782
rect 11670 3780 11726 3782
rect 11750 3780 11806 3782
rect 15212 3834 15268 3836
rect 15292 3834 15348 3836
rect 15372 3834 15428 3836
rect 15452 3834 15508 3836
rect 15212 3782 15258 3834
rect 15258 3782 15268 3834
rect 15292 3782 15322 3834
rect 15322 3782 15334 3834
rect 15334 3782 15348 3834
rect 15372 3782 15386 3834
rect 15386 3782 15398 3834
rect 15398 3782 15428 3834
rect 15452 3782 15462 3834
rect 15462 3782 15508 3834
rect 15212 3780 15268 3782
rect 15292 3780 15348 3782
rect 15372 3780 15428 3782
rect 15452 3780 15508 3782
rect 9659 3290 9715 3292
rect 9739 3290 9795 3292
rect 9819 3290 9875 3292
rect 9899 3290 9955 3292
rect 9659 3238 9705 3290
rect 9705 3238 9715 3290
rect 9739 3238 9769 3290
rect 9769 3238 9781 3290
rect 9781 3238 9795 3290
rect 9819 3238 9833 3290
rect 9833 3238 9845 3290
rect 9845 3238 9875 3290
rect 9899 3238 9909 3290
rect 9909 3238 9955 3290
rect 9659 3236 9715 3238
rect 9739 3236 9795 3238
rect 9819 3236 9875 3238
rect 9899 3236 9955 3238
rect 13361 3290 13417 3292
rect 13441 3290 13497 3292
rect 13521 3290 13577 3292
rect 13601 3290 13657 3292
rect 13361 3238 13407 3290
rect 13407 3238 13417 3290
rect 13441 3238 13471 3290
rect 13471 3238 13483 3290
rect 13483 3238 13497 3290
rect 13521 3238 13535 3290
rect 13535 3238 13547 3290
rect 13547 3238 13577 3290
rect 13601 3238 13611 3290
rect 13611 3238 13657 3290
rect 13361 3236 13417 3238
rect 13441 3236 13497 3238
rect 13521 3236 13577 3238
rect 13601 3236 13657 3238
rect 4106 2746 4162 2748
rect 4186 2746 4242 2748
rect 4266 2746 4322 2748
rect 4346 2746 4402 2748
rect 4106 2694 4152 2746
rect 4152 2694 4162 2746
rect 4186 2694 4216 2746
rect 4216 2694 4228 2746
rect 4228 2694 4242 2746
rect 4266 2694 4280 2746
rect 4280 2694 4292 2746
rect 4292 2694 4322 2746
rect 4346 2694 4356 2746
rect 4356 2694 4402 2746
rect 4106 2692 4162 2694
rect 4186 2692 4242 2694
rect 4266 2692 4322 2694
rect 4346 2692 4402 2694
rect 7808 2746 7864 2748
rect 7888 2746 7944 2748
rect 7968 2746 8024 2748
rect 8048 2746 8104 2748
rect 7808 2694 7854 2746
rect 7854 2694 7864 2746
rect 7888 2694 7918 2746
rect 7918 2694 7930 2746
rect 7930 2694 7944 2746
rect 7968 2694 7982 2746
rect 7982 2694 7994 2746
rect 7994 2694 8024 2746
rect 8048 2694 8058 2746
rect 8058 2694 8104 2746
rect 7808 2692 7864 2694
rect 7888 2692 7944 2694
rect 7968 2692 8024 2694
rect 8048 2692 8104 2694
rect 11510 2746 11566 2748
rect 11590 2746 11646 2748
rect 11670 2746 11726 2748
rect 11750 2746 11806 2748
rect 2255 2202 2311 2204
rect 2335 2202 2391 2204
rect 2415 2202 2471 2204
rect 2495 2202 2551 2204
rect 2255 2150 2301 2202
rect 2301 2150 2311 2202
rect 2335 2150 2365 2202
rect 2365 2150 2377 2202
rect 2377 2150 2391 2202
rect 2415 2150 2429 2202
rect 2429 2150 2441 2202
rect 2441 2150 2471 2202
rect 2495 2150 2505 2202
rect 2505 2150 2551 2202
rect 2255 2148 2311 2150
rect 2335 2148 2391 2150
rect 2415 2148 2471 2150
rect 2495 2148 2551 2150
rect 5957 2202 6013 2204
rect 6037 2202 6093 2204
rect 6117 2202 6173 2204
rect 6197 2202 6253 2204
rect 5957 2150 6003 2202
rect 6003 2150 6013 2202
rect 6037 2150 6067 2202
rect 6067 2150 6079 2202
rect 6079 2150 6093 2202
rect 6117 2150 6131 2202
rect 6131 2150 6143 2202
rect 6143 2150 6173 2202
rect 6197 2150 6207 2202
rect 6207 2150 6253 2202
rect 5957 2148 6013 2150
rect 6037 2148 6093 2150
rect 6117 2148 6173 2150
rect 6197 2148 6253 2150
rect 4106 1658 4162 1660
rect 4186 1658 4242 1660
rect 4266 1658 4322 1660
rect 4346 1658 4402 1660
rect 4106 1606 4152 1658
rect 4152 1606 4162 1658
rect 4186 1606 4216 1658
rect 4216 1606 4228 1658
rect 4228 1606 4242 1658
rect 4266 1606 4280 1658
rect 4280 1606 4292 1658
rect 4292 1606 4322 1658
rect 4346 1606 4356 1658
rect 4356 1606 4402 1658
rect 4106 1604 4162 1606
rect 4186 1604 4242 1606
rect 4266 1604 4322 1606
rect 4346 1604 4402 1606
rect 7808 1658 7864 1660
rect 7888 1658 7944 1660
rect 7968 1658 8024 1660
rect 8048 1658 8104 1660
rect 7808 1606 7854 1658
rect 7854 1606 7864 1658
rect 7888 1606 7918 1658
rect 7918 1606 7930 1658
rect 7930 1606 7944 1658
rect 7968 1606 7982 1658
rect 7982 1606 7994 1658
rect 7994 1606 8024 1658
rect 8048 1606 8058 1658
rect 8058 1606 8104 1658
rect 7808 1604 7864 1606
rect 7888 1604 7944 1606
rect 7968 1604 8024 1606
rect 8048 1604 8104 1606
rect 2255 1114 2311 1116
rect 2335 1114 2391 1116
rect 2415 1114 2471 1116
rect 2495 1114 2551 1116
rect 2255 1062 2301 1114
rect 2301 1062 2311 1114
rect 2335 1062 2365 1114
rect 2365 1062 2377 1114
rect 2377 1062 2391 1114
rect 2415 1062 2429 1114
rect 2429 1062 2441 1114
rect 2441 1062 2471 1114
rect 2495 1062 2505 1114
rect 2505 1062 2551 1114
rect 2255 1060 2311 1062
rect 2335 1060 2391 1062
rect 2415 1060 2471 1062
rect 2495 1060 2551 1062
rect 5957 1114 6013 1116
rect 6037 1114 6093 1116
rect 6117 1114 6173 1116
rect 6197 1114 6253 1116
rect 5957 1062 6003 1114
rect 6003 1062 6013 1114
rect 6037 1062 6067 1114
rect 6067 1062 6079 1114
rect 6079 1062 6093 1114
rect 6117 1062 6131 1114
rect 6131 1062 6143 1114
rect 6143 1062 6173 1114
rect 6197 1062 6207 1114
rect 6207 1062 6253 1114
rect 5957 1060 6013 1062
rect 6037 1060 6093 1062
rect 6117 1060 6173 1062
rect 6197 1060 6253 1062
rect 11510 2694 11556 2746
rect 11556 2694 11566 2746
rect 11590 2694 11620 2746
rect 11620 2694 11632 2746
rect 11632 2694 11646 2746
rect 11670 2694 11684 2746
rect 11684 2694 11696 2746
rect 11696 2694 11726 2746
rect 11750 2694 11760 2746
rect 11760 2694 11806 2746
rect 11510 2692 11566 2694
rect 11590 2692 11646 2694
rect 11670 2692 11726 2694
rect 11750 2692 11806 2694
rect 15212 2746 15268 2748
rect 15292 2746 15348 2748
rect 15372 2746 15428 2748
rect 15452 2746 15508 2748
rect 15212 2694 15258 2746
rect 15258 2694 15268 2746
rect 15292 2694 15322 2746
rect 15322 2694 15334 2746
rect 15334 2694 15348 2746
rect 15372 2694 15386 2746
rect 15386 2694 15398 2746
rect 15398 2694 15428 2746
rect 15452 2694 15462 2746
rect 15462 2694 15508 2746
rect 15212 2692 15268 2694
rect 15292 2692 15348 2694
rect 15372 2692 15428 2694
rect 15452 2692 15508 2694
rect 9659 2202 9715 2204
rect 9739 2202 9795 2204
rect 9819 2202 9875 2204
rect 9899 2202 9955 2204
rect 9659 2150 9705 2202
rect 9705 2150 9715 2202
rect 9739 2150 9769 2202
rect 9769 2150 9781 2202
rect 9781 2150 9795 2202
rect 9819 2150 9833 2202
rect 9833 2150 9845 2202
rect 9845 2150 9875 2202
rect 9899 2150 9909 2202
rect 9909 2150 9955 2202
rect 9659 2148 9715 2150
rect 9739 2148 9795 2150
rect 9819 2148 9875 2150
rect 9899 2148 9955 2150
rect 13361 2202 13417 2204
rect 13441 2202 13497 2204
rect 13521 2202 13577 2204
rect 13601 2202 13657 2204
rect 13361 2150 13407 2202
rect 13407 2150 13417 2202
rect 13441 2150 13471 2202
rect 13471 2150 13483 2202
rect 13483 2150 13497 2202
rect 13521 2150 13535 2202
rect 13535 2150 13547 2202
rect 13547 2150 13577 2202
rect 13601 2150 13611 2202
rect 13611 2150 13657 2202
rect 13361 2148 13417 2150
rect 13441 2148 13497 2150
rect 13521 2148 13577 2150
rect 13601 2148 13657 2150
rect 11510 1658 11566 1660
rect 11590 1658 11646 1660
rect 11670 1658 11726 1660
rect 11750 1658 11806 1660
rect 11510 1606 11556 1658
rect 11556 1606 11566 1658
rect 11590 1606 11620 1658
rect 11620 1606 11632 1658
rect 11632 1606 11646 1658
rect 11670 1606 11684 1658
rect 11684 1606 11696 1658
rect 11696 1606 11726 1658
rect 11750 1606 11760 1658
rect 11760 1606 11806 1658
rect 11510 1604 11566 1606
rect 11590 1604 11646 1606
rect 11670 1604 11726 1606
rect 11750 1604 11806 1606
rect 15212 1658 15268 1660
rect 15292 1658 15348 1660
rect 15372 1658 15428 1660
rect 15452 1658 15508 1660
rect 15212 1606 15258 1658
rect 15258 1606 15268 1658
rect 15292 1606 15322 1658
rect 15322 1606 15334 1658
rect 15334 1606 15348 1658
rect 15372 1606 15386 1658
rect 15386 1606 15398 1658
rect 15398 1606 15428 1658
rect 15452 1606 15462 1658
rect 15462 1606 15508 1658
rect 15212 1604 15268 1606
rect 15292 1604 15348 1606
rect 15372 1604 15428 1606
rect 15452 1604 15508 1606
rect 9659 1114 9715 1116
rect 9739 1114 9795 1116
rect 9819 1114 9875 1116
rect 9899 1114 9955 1116
rect 9659 1062 9705 1114
rect 9705 1062 9715 1114
rect 9739 1062 9769 1114
rect 9769 1062 9781 1114
rect 9781 1062 9795 1114
rect 9819 1062 9833 1114
rect 9833 1062 9845 1114
rect 9845 1062 9875 1114
rect 9899 1062 9909 1114
rect 9909 1062 9955 1114
rect 9659 1060 9715 1062
rect 9739 1060 9795 1062
rect 9819 1060 9875 1062
rect 9899 1060 9955 1062
rect 13361 1114 13417 1116
rect 13441 1114 13497 1116
rect 13521 1114 13577 1116
rect 13601 1114 13657 1116
rect 13361 1062 13407 1114
rect 13407 1062 13417 1114
rect 13441 1062 13471 1114
rect 13471 1062 13483 1114
rect 13483 1062 13497 1114
rect 13521 1062 13535 1114
rect 13535 1062 13547 1114
rect 13547 1062 13577 1114
rect 13601 1062 13611 1114
rect 13611 1062 13657 1114
rect 13361 1060 13417 1062
rect 13441 1060 13497 1062
rect 13521 1060 13577 1062
rect 13601 1060 13657 1062
rect 4106 570 4162 572
rect 4186 570 4242 572
rect 4266 570 4322 572
rect 4346 570 4402 572
rect 4106 518 4152 570
rect 4152 518 4162 570
rect 4186 518 4216 570
rect 4216 518 4228 570
rect 4228 518 4242 570
rect 4266 518 4280 570
rect 4280 518 4292 570
rect 4292 518 4322 570
rect 4346 518 4356 570
rect 4356 518 4402 570
rect 4106 516 4162 518
rect 4186 516 4242 518
rect 4266 516 4322 518
rect 4346 516 4402 518
rect 7808 570 7864 572
rect 7888 570 7944 572
rect 7968 570 8024 572
rect 8048 570 8104 572
rect 7808 518 7854 570
rect 7854 518 7864 570
rect 7888 518 7918 570
rect 7918 518 7930 570
rect 7930 518 7944 570
rect 7968 518 7982 570
rect 7982 518 7994 570
rect 7994 518 8024 570
rect 8048 518 8058 570
rect 8058 518 8104 570
rect 7808 516 7864 518
rect 7888 516 7944 518
rect 7968 516 8024 518
rect 8048 516 8104 518
rect 11510 570 11566 572
rect 11590 570 11646 572
rect 11670 570 11726 572
rect 11750 570 11806 572
rect 11510 518 11556 570
rect 11556 518 11566 570
rect 11590 518 11620 570
rect 11620 518 11632 570
rect 11632 518 11646 570
rect 11670 518 11684 570
rect 11684 518 11696 570
rect 11696 518 11726 570
rect 11750 518 11760 570
rect 11760 518 11806 570
rect 11510 516 11566 518
rect 11590 516 11646 518
rect 11670 516 11726 518
rect 11750 516 11806 518
rect 15212 570 15268 572
rect 15292 570 15348 572
rect 15372 570 15428 572
rect 15452 570 15508 572
rect 15212 518 15258 570
rect 15258 518 15268 570
rect 15292 518 15322 570
rect 15322 518 15334 570
rect 15334 518 15348 570
rect 15372 518 15386 570
rect 15386 518 15398 570
rect 15398 518 15428 570
rect 15452 518 15462 570
rect 15462 518 15508 570
rect 15212 516 15268 518
rect 15292 516 15348 518
rect 15372 516 15428 518
rect 15452 516 15508 518
<< metal3 >>
rect 2245 15264 2561 15265
rect 2245 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2561 15264
rect 2245 15199 2561 15200
rect 5947 15264 6263 15265
rect 5947 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6263 15264
rect 5947 15199 6263 15200
rect 9649 15264 9965 15265
rect 9649 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9965 15264
rect 9649 15199 9965 15200
rect 13351 15264 13667 15265
rect 13351 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13667 15264
rect 13351 15199 13667 15200
rect 4096 14720 4412 14721
rect 4096 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4412 14720
rect 4096 14655 4412 14656
rect 7798 14720 8114 14721
rect 7798 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8114 14720
rect 7798 14655 8114 14656
rect 11500 14720 11816 14721
rect 11500 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11816 14720
rect 11500 14655 11816 14656
rect 15202 14720 15518 14721
rect 15202 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15518 14720
rect 15202 14655 15518 14656
rect 2245 14176 2561 14177
rect 2245 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2561 14176
rect 2245 14111 2561 14112
rect 5947 14176 6263 14177
rect 5947 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6263 14176
rect 5947 14111 6263 14112
rect 9649 14176 9965 14177
rect 9649 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9965 14176
rect 9649 14111 9965 14112
rect 13351 14176 13667 14177
rect 13351 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13667 14176
rect 13351 14111 13667 14112
rect 4096 13632 4412 13633
rect 4096 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4412 13632
rect 4096 13567 4412 13568
rect 7798 13632 8114 13633
rect 7798 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8114 13632
rect 7798 13567 8114 13568
rect 11500 13632 11816 13633
rect 11500 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11816 13632
rect 11500 13567 11816 13568
rect 15202 13632 15518 13633
rect 15202 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15518 13632
rect 15202 13567 15518 13568
rect 2245 13088 2561 13089
rect 2245 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2561 13088
rect 2245 13023 2561 13024
rect 5947 13088 6263 13089
rect 5947 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6263 13088
rect 5947 13023 6263 13024
rect 9649 13088 9965 13089
rect 9649 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9965 13088
rect 9649 13023 9965 13024
rect 13351 13088 13667 13089
rect 13351 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13667 13088
rect 13351 13023 13667 13024
rect 4096 12544 4412 12545
rect 4096 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4412 12544
rect 4096 12479 4412 12480
rect 7798 12544 8114 12545
rect 7798 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8114 12544
rect 7798 12479 8114 12480
rect 11500 12544 11816 12545
rect 11500 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11816 12544
rect 11500 12479 11816 12480
rect 15202 12544 15518 12545
rect 15202 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15518 12544
rect 15202 12479 15518 12480
rect 6453 12474 6519 12477
rect 6318 12472 6519 12474
rect 6318 12416 6458 12472
rect 6514 12416 6519 12472
rect 6318 12414 6519 12416
rect 2681 12338 2747 12341
rect 6318 12338 6378 12414
rect 6453 12411 6519 12414
rect 2681 12336 6378 12338
rect 2681 12280 2686 12336
rect 2742 12280 6378 12336
rect 2681 12278 6378 12280
rect 2681 12275 2747 12278
rect 2245 12000 2561 12001
rect 2245 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2561 12000
rect 2245 11935 2561 11936
rect 5947 12000 6263 12001
rect 5947 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6263 12000
rect 5947 11935 6263 11936
rect 9649 12000 9965 12001
rect 9649 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9965 12000
rect 9649 11935 9965 11936
rect 13351 12000 13667 12001
rect 13351 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13667 12000
rect 13351 11935 13667 11936
rect 4096 11456 4412 11457
rect 4096 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4412 11456
rect 4096 11391 4412 11392
rect 7798 11456 8114 11457
rect 7798 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8114 11456
rect 7798 11391 8114 11392
rect 11500 11456 11816 11457
rect 11500 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11816 11456
rect 11500 11391 11816 11392
rect 15202 11456 15518 11457
rect 15202 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15518 11456
rect 15202 11391 15518 11392
rect 2245 10912 2561 10913
rect 2245 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2561 10912
rect 2245 10847 2561 10848
rect 5947 10912 6263 10913
rect 5947 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6263 10912
rect 5947 10847 6263 10848
rect 9649 10912 9965 10913
rect 9649 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9965 10912
rect 9649 10847 9965 10848
rect 13351 10912 13667 10913
rect 13351 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13667 10912
rect 13351 10847 13667 10848
rect 4096 10368 4412 10369
rect 4096 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4412 10368
rect 4096 10303 4412 10304
rect 7798 10368 8114 10369
rect 7798 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8114 10368
rect 7798 10303 8114 10304
rect 11500 10368 11816 10369
rect 11500 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11816 10368
rect 11500 10303 11816 10304
rect 15202 10368 15518 10369
rect 15202 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15518 10368
rect 15202 10303 15518 10304
rect 2245 9824 2561 9825
rect 2245 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2561 9824
rect 2245 9759 2561 9760
rect 5947 9824 6263 9825
rect 5947 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6263 9824
rect 5947 9759 6263 9760
rect 9649 9824 9965 9825
rect 9649 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9965 9824
rect 9649 9759 9965 9760
rect 13351 9824 13667 9825
rect 13351 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13667 9824
rect 13351 9759 13667 9760
rect 4096 9280 4412 9281
rect 4096 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4412 9280
rect 4096 9215 4412 9216
rect 7798 9280 8114 9281
rect 7798 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8114 9280
rect 7798 9215 8114 9216
rect 11500 9280 11816 9281
rect 11500 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11816 9280
rect 11500 9215 11816 9216
rect 15202 9280 15518 9281
rect 15202 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15518 9280
rect 15202 9215 15518 9216
rect 2245 8736 2561 8737
rect 2245 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2561 8736
rect 2245 8671 2561 8672
rect 5947 8736 6263 8737
rect 5947 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6263 8736
rect 5947 8671 6263 8672
rect 9649 8736 9965 8737
rect 9649 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9965 8736
rect 9649 8671 9965 8672
rect 13351 8736 13667 8737
rect 13351 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13667 8736
rect 13351 8671 13667 8672
rect 4096 8192 4412 8193
rect 4096 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4412 8192
rect 4096 8127 4412 8128
rect 7798 8192 8114 8193
rect 7798 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8114 8192
rect 7798 8127 8114 8128
rect 11500 8192 11816 8193
rect 11500 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11816 8192
rect 11500 8127 11816 8128
rect 15202 8192 15518 8193
rect 15202 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15518 8192
rect 15202 8127 15518 8128
rect 2245 7648 2561 7649
rect 2245 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2561 7648
rect 2245 7583 2561 7584
rect 5947 7648 6263 7649
rect 5947 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6263 7648
rect 5947 7583 6263 7584
rect 9649 7648 9965 7649
rect 9649 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9965 7648
rect 9649 7583 9965 7584
rect 13351 7648 13667 7649
rect 13351 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13667 7648
rect 13351 7583 13667 7584
rect 4096 7104 4412 7105
rect 4096 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4412 7104
rect 4096 7039 4412 7040
rect 7798 7104 8114 7105
rect 7798 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8114 7104
rect 7798 7039 8114 7040
rect 11500 7104 11816 7105
rect 11500 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11816 7104
rect 11500 7039 11816 7040
rect 15202 7104 15518 7105
rect 15202 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15518 7104
rect 15202 7039 15518 7040
rect 2245 6560 2561 6561
rect 2245 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2561 6560
rect 2245 6495 2561 6496
rect 5947 6560 6263 6561
rect 5947 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6263 6560
rect 5947 6495 6263 6496
rect 9649 6560 9965 6561
rect 9649 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9965 6560
rect 9649 6495 9965 6496
rect 13351 6560 13667 6561
rect 13351 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13667 6560
rect 13351 6495 13667 6496
rect 4096 6016 4412 6017
rect 4096 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4412 6016
rect 4096 5951 4412 5952
rect 7798 6016 8114 6017
rect 7798 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8114 6016
rect 7798 5951 8114 5952
rect 11500 6016 11816 6017
rect 11500 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11816 6016
rect 11500 5951 11816 5952
rect 15202 6016 15518 6017
rect 15202 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15518 6016
rect 15202 5951 15518 5952
rect 2245 5472 2561 5473
rect 2245 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2561 5472
rect 2245 5407 2561 5408
rect 5947 5472 6263 5473
rect 5947 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6263 5472
rect 5947 5407 6263 5408
rect 9649 5472 9965 5473
rect 9649 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9965 5472
rect 9649 5407 9965 5408
rect 13351 5472 13667 5473
rect 13351 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13667 5472
rect 13351 5407 13667 5408
rect 4096 4928 4412 4929
rect 4096 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4412 4928
rect 4096 4863 4412 4864
rect 7798 4928 8114 4929
rect 7798 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8114 4928
rect 7798 4863 8114 4864
rect 11500 4928 11816 4929
rect 11500 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11816 4928
rect 11500 4863 11816 4864
rect 15202 4928 15518 4929
rect 15202 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15518 4928
rect 15202 4863 15518 4864
rect 2245 4384 2561 4385
rect 2245 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2561 4384
rect 2245 4319 2561 4320
rect 5947 4384 6263 4385
rect 5947 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6263 4384
rect 5947 4319 6263 4320
rect 9649 4384 9965 4385
rect 9649 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9965 4384
rect 9649 4319 9965 4320
rect 13351 4384 13667 4385
rect 13351 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13667 4384
rect 13351 4319 13667 4320
rect 4096 3840 4412 3841
rect 4096 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4412 3840
rect 4096 3775 4412 3776
rect 7798 3840 8114 3841
rect 7798 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8114 3840
rect 7798 3775 8114 3776
rect 11500 3840 11816 3841
rect 11500 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11816 3840
rect 11500 3775 11816 3776
rect 15202 3840 15518 3841
rect 15202 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15518 3840
rect 15202 3775 15518 3776
rect 2245 3296 2561 3297
rect 2245 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2561 3296
rect 2245 3231 2561 3232
rect 5947 3296 6263 3297
rect 5947 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6263 3296
rect 5947 3231 6263 3232
rect 9649 3296 9965 3297
rect 9649 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9965 3296
rect 9649 3231 9965 3232
rect 13351 3296 13667 3297
rect 13351 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13667 3296
rect 13351 3231 13667 3232
rect 4096 2752 4412 2753
rect 4096 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4412 2752
rect 4096 2687 4412 2688
rect 7798 2752 8114 2753
rect 7798 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8114 2752
rect 7798 2687 8114 2688
rect 11500 2752 11816 2753
rect 11500 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11816 2752
rect 11500 2687 11816 2688
rect 15202 2752 15518 2753
rect 15202 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15518 2752
rect 15202 2687 15518 2688
rect 2245 2208 2561 2209
rect 2245 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2561 2208
rect 2245 2143 2561 2144
rect 5947 2208 6263 2209
rect 5947 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6263 2208
rect 5947 2143 6263 2144
rect 9649 2208 9965 2209
rect 9649 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9965 2208
rect 9649 2143 9965 2144
rect 13351 2208 13667 2209
rect 13351 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13667 2208
rect 13351 2143 13667 2144
rect 4096 1664 4412 1665
rect 4096 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4412 1664
rect 4096 1599 4412 1600
rect 7798 1664 8114 1665
rect 7798 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8114 1664
rect 7798 1599 8114 1600
rect 11500 1664 11816 1665
rect 11500 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11816 1664
rect 11500 1599 11816 1600
rect 15202 1664 15518 1665
rect 15202 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15518 1664
rect 15202 1599 15518 1600
rect 2245 1120 2561 1121
rect 2245 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2561 1120
rect 2245 1055 2561 1056
rect 5947 1120 6263 1121
rect 5947 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6263 1120
rect 5947 1055 6263 1056
rect 9649 1120 9965 1121
rect 9649 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9965 1120
rect 9649 1055 9965 1056
rect 13351 1120 13667 1121
rect 13351 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13667 1120
rect 13351 1055 13667 1056
rect 4096 576 4412 577
rect 4096 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4412 576
rect 4096 511 4412 512
rect 7798 576 8114 577
rect 7798 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8114 576
rect 7798 511 8114 512
rect 11500 576 11816 577
rect 11500 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11816 576
rect 11500 511 11816 512
rect 15202 576 15518 577
rect 15202 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15518 576
rect 15202 511 15518 512
<< via3 >>
rect 2251 15260 2315 15264
rect 2251 15204 2255 15260
rect 2255 15204 2311 15260
rect 2311 15204 2315 15260
rect 2251 15200 2315 15204
rect 2331 15260 2395 15264
rect 2331 15204 2335 15260
rect 2335 15204 2391 15260
rect 2391 15204 2395 15260
rect 2331 15200 2395 15204
rect 2411 15260 2475 15264
rect 2411 15204 2415 15260
rect 2415 15204 2471 15260
rect 2471 15204 2475 15260
rect 2411 15200 2475 15204
rect 2491 15260 2555 15264
rect 2491 15204 2495 15260
rect 2495 15204 2551 15260
rect 2551 15204 2555 15260
rect 2491 15200 2555 15204
rect 5953 15260 6017 15264
rect 5953 15204 5957 15260
rect 5957 15204 6013 15260
rect 6013 15204 6017 15260
rect 5953 15200 6017 15204
rect 6033 15260 6097 15264
rect 6033 15204 6037 15260
rect 6037 15204 6093 15260
rect 6093 15204 6097 15260
rect 6033 15200 6097 15204
rect 6113 15260 6177 15264
rect 6113 15204 6117 15260
rect 6117 15204 6173 15260
rect 6173 15204 6177 15260
rect 6113 15200 6177 15204
rect 6193 15260 6257 15264
rect 6193 15204 6197 15260
rect 6197 15204 6253 15260
rect 6253 15204 6257 15260
rect 6193 15200 6257 15204
rect 9655 15260 9719 15264
rect 9655 15204 9659 15260
rect 9659 15204 9715 15260
rect 9715 15204 9719 15260
rect 9655 15200 9719 15204
rect 9735 15260 9799 15264
rect 9735 15204 9739 15260
rect 9739 15204 9795 15260
rect 9795 15204 9799 15260
rect 9735 15200 9799 15204
rect 9815 15260 9879 15264
rect 9815 15204 9819 15260
rect 9819 15204 9875 15260
rect 9875 15204 9879 15260
rect 9815 15200 9879 15204
rect 9895 15260 9959 15264
rect 9895 15204 9899 15260
rect 9899 15204 9955 15260
rect 9955 15204 9959 15260
rect 9895 15200 9959 15204
rect 13357 15260 13421 15264
rect 13357 15204 13361 15260
rect 13361 15204 13417 15260
rect 13417 15204 13421 15260
rect 13357 15200 13421 15204
rect 13437 15260 13501 15264
rect 13437 15204 13441 15260
rect 13441 15204 13497 15260
rect 13497 15204 13501 15260
rect 13437 15200 13501 15204
rect 13517 15260 13581 15264
rect 13517 15204 13521 15260
rect 13521 15204 13577 15260
rect 13577 15204 13581 15260
rect 13517 15200 13581 15204
rect 13597 15260 13661 15264
rect 13597 15204 13601 15260
rect 13601 15204 13657 15260
rect 13657 15204 13661 15260
rect 13597 15200 13661 15204
rect 4102 14716 4166 14720
rect 4102 14660 4106 14716
rect 4106 14660 4162 14716
rect 4162 14660 4166 14716
rect 4102 14656 4166 14660
rect 4182 14716 4246 14720
rect 4182 14660 4186 14716
rect 4186 14660 4242 14716
rect 4242 14660 4246 14716
rect 4182 14656 4246 14660
rect 4262 14716 4326 14720
rect 4262 14660 4266 14716
rect 4266 14660 4322 14716
rect 4322 14660 4326 14716
rect 4262 14656 4326 14660
rect 4342 14716 4406 14720
rect 4342 14660 4346 14716
rect 4346 14660 4402 14716
rect 4402 14660 4406 14716
rect 4342 14656 4406 14660
rect 7804 14716 7868 14720
rect 7804 14660 7808 14716
rect 7808 14660 7864 14716
rect 7864 14660 7868 14716
rect 7804 14656 7868 14660
rect 7884 14716 7948 14720
rect 7884 14660 7888 14716
rect 7888 14660 7944 14716
rect 7944 14660 7948 14716
rect 7884 14656 7948 14660
rect 7964 14716 8028 14720
rect 7964 14660 7968 14716
rect 7968 14660 8024 14716
rect 8024 14660 8028 14716
rect 7964 14656 8028 14660
rect 8044 14716 8108 14720
rect 8044 14660 8048 14716
rect 8048 14660 8104 14716
rect 8104 14660 8108 14716
rect 8044 14656 8108 14660
rect 11506 14716 11570 14720
rect 11506 14660 11510 14716
rect 11510 14660 11566 14716
rect 11566 14660 11570 14716
rect 11506 14656 11570 14660
rect 11586 14716 11650 14720
rect 11586 14660 11590 14716
rect 11590 14660 11646 14716
rect 11646 14660 11650 14716
rect 11586 14656 11650 14660
rect 11666 14716 11730 14720
rect 11666 14660 11670 14716
rect 11670 14660 11726 14716
rect 11726 14660 11730 14716
rect 11666 14656 11730 14660
rect 11746 14716 11810 14720
rect 11746 14660 11750 14716
rect 11750 14660 11806 14716
rect 11806 14660 11810 14716
rect 11746 14656 11810 14660
rect 15208 14716 15272 14720
rect 15208 14660 15212 14716
rect 15212 14660 15268 14716
rect 15268 14660 15272 14716
rect 15208 14656 15272 14660
rect 15288 14716 15352 14720
rect 15288 14660 15292 14716
rect 15292 14660 15348 14716
rect 15348 14660 15352 14716
rect 15288 14656 15352 14660
rect 15368 14716 15432 14720
rect 15368 14660 15372 14716
rect 15372 14660 15428 14716
rect 15428 14660 15432 14716
rect 15368 14656 15432 14660
rect 15448 14716 15512 14720
rect 15448 14660 15452 14716
rect 15452 14660 15508 14716
rect 15508 14660 15512 14716
rect 15448 14656 15512 14660
rect 2251 14172 2315 14176
rect 2251 14116 2255 14172
rect 2255 14116 2311 14172
rect 2311 14116 2315 14172
rect 2251 14112 2315 14116
rect 2331 14172 2395 14176
rect 2331 14116 2335 14172
rect 2335 14116 2391 14172
rect 2391 14116 2395 14172
rect 2331 14112 2395 14116
rect 2411 14172 2475 14176
rect 2411 14116 2415 14172
rect 2415 14116 2471 14172
rect 2471 14116 2475 14172
rect 2411 14112 2475 14116
rect 2491 14172 2555 14176
rect 2491 14116 2495 14172
rect 2495 14116 2551 14172
rect 2551 14116 2555 14172
rect 2491 14112 2555 14116
rect 5953 14172 6017 14176
rect 5953 14116 5957 14172
rect 5957 14116 6013 14172
rect 6013 14116 6017 14172
rect 5953 14112 6017 14116
rect 6033 14172 6097 14176
rect 6033 14116 6037 14172
rect 6037 14116 6093 14172
rect 6093 14116 6097 14172
rect 6033 14112 6097 14116
rect 6113 14172 6177 14176
rect 6113 14116 6117 14172
rect 6117 14116 6173 14172
rect 6173 14116 6177 14172
rect 6113 14112 6177 14116
rect 6193 14172 6257 14176
rect 6193 14116 6197 14172
rect 6197 14116 6253 14172
rect 6253 14116 6257 14172
rect 6193 14112 6257 14116
rect 9655 14172 9719 14176
rect 9655 14116 9659 14172
rect 9659 14116 9715 14172
rect 9715 14116 9719 14172
rect 9655 14112 9719 14116
rect 9735 14172 9799 14176
rect 9735 14116 9739 14172
rect 9739 14116 9795 14172
rect 9795 14116 9799 14172
rect 9735 14112 9799 14116
rect 9815 14172 9879 14176
rect 9815 14116 9819 14172
rect 9819 14116 9875 14172
rect 9875 14116 9879 14172
rect 9815 14112 9879 14116
rect 9895 14172 9959 14176
rect 9895 14116 9899 14172
rect 9899 14116 9955 14172
rect 9955 14116 9959 14172
rect 9895 14112 9959 14116
rect 13357 14172 13421 14176
rect 13357 14116 13361 14172
rect 13361 14116 13417 14172
rect 13417 14116 13421 14172
rect 13357 14112 13421 14116
rect 13437 14172 13501 14176
rect 13437 14116 13441 14172
rect 13441 14116 13497 14172
rect 13497 14116 13501 14172
rect 13437 14112 13501 14116
rect 13517 14172 13581 14176
rect 13517 14116 13521 14172
rect 13521 14116 13577 14172
rect 13577 14116 13581 14172
rect 13517 14112 13581 14116
rect 13597 14172 13661 14176
rect 13597 14116 13601 14172
rect 13601 14116 13657 14172
rect 13657 14116 13661 14172
rect 13597 14112 13661 14116
rect 4102 13628 4166 13632
rect 4102 13572 4106 13628
rect 4106 13572 4162 13628
rect 4162 13572 4166 13628
rect 4102 13568 4166 13572
rect 4182 13628 4246 13632
rect 4182 13572 4186 13628
rect 4186 13572 4242 13628
rect 4242 13572 4246 13628
rect 4182 13568 4246 13572
rect 4262 13628 4326 13632
rect 4262 13572 4266 13628
rect 4266 13572 4322 13628
rect 4322 13572 4326 13628
rect 4262 13568 4326 13572
rect 4342 13628 4406 13632
rect 4342 13572 4346 13628
rect 4346 13572 4402 13628
rect 4402 13572 4406 13628
rect 4342 13568 4406 13572
rect 7804 13628 7868 13632
rect 7804 13572 7808 13628
rect 7808 13572 7864 13628
rect 7864 13572 7868 13628
rect 7804 13568 7868 13572
rect 7884 13628 7948 13632
rect 7884 13572 7888 13628
rect 7888 13572 7944 13628
rect 7944 13572 7948 13628
rect 7884 13568 7948 13572
rect 7964 13628 8028 13632
rect 7964 13572 7968 13628
rect 7968 13572 8024 13628
rect 8024 13572 8028 13628
rect 7964 13568 8028 13572
rect 8044 13628 8108 13632
rect 8044 13572 8048 13628
rect 8048 13572 8104 13628
rect 8104 13572 8108 13628
rect 8044 13568 8108 13572
rect 11506 13628 11570 13632
rect 11506 13572 11510 13628
rect 11510 13572 11566 13628
rect 11566 13572 11570 13628
rect 11506 13568 11570 13572
rect 11586 13628 11650 13632
rect 11586 13572 11590 13628
rect 11590 13572 11646 13628
rect 11646 13572 11650 13628
rect 11586 13568 11650 13572
rect 11666 13628 11730 13632
rect 11666 13572 11670 13628
rect 11670 13572 11726 13628
rect 11726 13572 11730 13628
rect 11666 13568 11730 13572
rect 11746 13628 11810 13632
rect 11746 13572 11750 13628
rect 11750 13572 11806 13628
rect 11806 13572 11810 13628
rect 11746 13568 11810 13572
rect 15208 13628 15272 13632
rect 15208 13572 15212 13628
rect 15212 13572 15268 13628
rect 15268 13572 15272 13628
rect 15208 13568 15272 13572
rect 15288 13628 15352 13632
rect 15288 13572 15292 13628
rect 15292 13572 15348 13628
rect 15348 13572 15352 13628
rect 15288 13568 15352 13572
rect 15368 13628 15432 13632
rect 15368 13572 15372 13628
rect 15372 13572 15428 13628
rect 15428 13572 15432 13628
rect 15368 13568 15432 13572
rect 15448 13628 15512 13632
rect 15448 13572 15452 13628
rect 15452 13572 15508 13628
rect 15508 13572 15512 13628
rect 15448 13568 15512 13572
rect 2251 13084 2315 13088
rect 2251 13028 2255 13084
rect 2255 13028 2311 13084
rect 2311 13028 2315 13084
rect 2251 13024 2315 13028
rect 2331 13084 2395 13088
rect 2331 13028 2335 13084
rect 2335 13028 2391 13084
rect 2391 13028 2395 13084
rect 2331 13024 2395 13028
rect 2411 13084 2475 13088
rect 2411 13028 2415 13084
rect 2415 13028 2471 13084
rect 2471 13028 2475 13084
rect 2411 13024 2475 13028
rect 2491 13084 2555 13088
rect 2491 13028 2495 13084
rect 2495 13028 2551 13084
rect 2551 13028 2555 13084
rect 2491 13024 2555 13028
rect 5953 13084 6017 13088
rect 5953 13028 5957 13084
rect 5957 13028 6013 13084
rect 6013 13028 6017 13084
rect 5953 13024 6017 13028
rect 6033 13084 6097 13088
rect 6033 13028 6037 13084
rect 6037 13028 6093 13084
rect 6093 13028 6097 13084
rect 6033 13024 6097 13028
rect 6113 13084 6177 13088
rect 6113 13028 6117 13084
rect 6117 13028 6173 13084
rect 6173 13028 6177 13084
rect 6113 13024 6177 13028
rect 6193 13084 6257 13088
rect 6193 13028 6197 13084
rect 6197 13028 6253 13084
rect 6253 13028 6257 13084
rect 6193 13024 6257 13028
rect 9655 13084 9719 13088
rect 9655 13028 9659 13084
rect 9659 13028 9715 13084
rect 9715 13028 9719 13084
rect 9655 13024 9719 13028
rect 9735 13084 9799 13088
rect 9735 13028 9739 13084
rect 9739 13028 9795 13084
rect 9795 13028 9799 13084
rect 9735 13024 9799 13028
rect 9815 13084 9879 13088
rect 9815 13028 9819 13084
rect 9819 13028 9875 13084
rect 9875 13028 9879 13084
rect 9815 13024 9879 13028
rect 9895 13084 9959 13088
rect 9895 13028 9899 13084
rect 9899 13028 9955 13084
rect 9955 13028 9959 13084
rect 9895 13024 9959 13028
rect 13357 13084 13421 13088
rect 13357 13028 13361 13084
rect 13361 13028 13417 13084
rect 13417 13028 13421 13084
rect 13357 13024 13421 13028
rect 13437 13084 13501 13088
rect 13437 13028 13441 13084
rect 13441 13028 13497 13084
rect 13497 13028 13501 13084
rect 13437 13024 13501 13028
rect 13517 13084 13581 13088
rect 13517 13028 13521 13084
rect 13521 13028 13577 13084
rect 13577 13028 13581 13084
rect 13517 13024 13581 13028
rect 13597 13084 13661 13088
rect 13597 13028 13601 13084
rect 13601 13028 13657 13084
rect 13657 13028 13661 13084
rect 13597 13024 13661 13028
rect 4102 12540 4166 12544
rect 4102 12484 4106 12540
rect 4106 12484 4162 12540
rect 4162 12484 4166 12540
rect 4102 12480 4166 12484
rect 4182 12540 4246 12544
rect 4182 12484 4186 12540
rect 4186 12484 4242 12540
rect 4242 12484 4246 12540
rect 4182 12480 4246 12484
rect 4262 12540 4326 12544
rect 4262 12484 4266 12540
rect 4266 12484 4322 12540
rect 4322 12484 4326 12540
rect 4262 12480 4326 12484
rect 4342 12540 4406 12544
rect 4342 12484 4346 12540
rect 4346 12484 4402 12540
rect 4402 12484 4406 12540
rect 4342 12480 4406 12484
rect 7804 12540 7868 12544
rect 7804 12484 7808 12540
rect 7808 12484 7864 12540
rect 7864 12484 7868 12540
rect 7804 12480 7868 12484
rect 7884 12540 7948 12544
rect 7884 12484 7888 12540
rect 7888 12484 7944 12540
rect 7944 12484 7948 12540
rect 7884 12480 7948 12484
rect 7964 12540 8028 12544
rect 7964 12484 7968 12540
rect 7968 12484 8024 12540
rect 8024 12484 8028 12540
rect 7964 12480 8028 12484
rect 8044 12540 8108 12544
rect 8044 12484 8048 12540
rect 8048 12484 8104 12540
rect 8104 12484 8108 12540
rect 8044 12480 8108 12484
rect 11506 12540 11570 12544
rect 11506 12484 11510 12540
rect 11510 12484 11566 12540
rect 11566 12484 11570 12540
rect 11506 12480 11570 12484
rect 11586 12540 11650 12544
rect 11586 12484 11590 12540
rect 11590 12484 11646 12540
rect 11646 12484 11650 12540
rect 11586 12480 11650 12484
rect 11666 12540 11730 12544
rect 11666 12484 11670 12540
rect 11670 12484 11726 12540
rect 11726 12484 11730 12540
rect 11666 12480 11730 12484
rect 11746 12540 11810 12544
rect 11746 12484 11750 12540
rect 11750 12484 11806 12540
rect 11806 12484 11810 12540
rect 11746 12480 11810 12484
rect 15208 12540 15272 12544
rect 15208 12484 15212 12540
rect 15212 12484 15268 12540
rect 15268 12484 15272 12540
rect 15208 12480 15272 12484
rect 15288 12540 15352 12544
rect 15288 12484 15292 12540
rect 15292 12484 15348 12540
rect 15348 12484 15352 12540
rect 15288 12480 15352 12484
rect 15368 12540 15432 12544
rect 15368 12484 15372 12540
rect 15372 12484 15428 12540
rect 15428 12484 15432 12540
rect 15368 12480 15432 12484
rect 15448 12540 15512 12544
rect 15448 12484 15452 12540
rect 15452 12484 15508 12540
rect 15508 12484 15512 12540
rect 15448 12480 15512 12484
rect 2251 11996 2315 12000
rect 2251 11940 2255 11996
rect 2255 11940 2311 11996
rect 2311 11940 2315 11996
rect 2251 11936 2315 11940
rect 2331 11996 2395 12000
rect 2331 11940 2335 11996
rect 2335 11940 2391 11996
rect 2391 11940 2395 11996
rect 2331 11936 2395 11940
rect 2411 11996 2475 12000
rect 2411 11940 2415 11996
rect 2415 11940 2471 11996
rect 2471 11940 2475 11996
rect 2411 11936 2475 11940
rect 2491 11996 2555 12000
rect 2491 11940 2495 11996
rect 2495 11940 2551 11996
rect 2551 11940 2555 11996
rect 2491 11936 2555 11940
rect 5953 11996 6017 12000
rect 5953 11940 5957 11996
rect 5957 11940 6013 11996
rect 6013 11940 6017 11996
rect 5953 11936 6017 11940
rect 6033 11996 6097 12000
rect 6033 11940 6037 11996
rect 6037 11940 6093 11996
rect 6093 11940 6097 11996
rect 6033 11936 6097 11940
rect 6113 11996 6177 12000
rect 6113 11940 6117 11996
rect 6117 11940 6173 11996
rect 6173 11940 6177 11996
rect 6113 11936 6177 11940
rect 6193 11996 6257 12000
rect 6193 11940 6197 11996
rect 6197 11940 6253 11996
rect 6253 11940 6257 11996
rect 6193 11936 6257 11940
rect 9655 11996 9719 12000
rect 9655 11940 9659 11996
rect 9659 11940 9715 11996
rect 9715 11940 9719 11996
rect 9655 11936 9719 11940
rect 9735 11996 9799 12000
rect 9735 11940 9739 11996
rect 9739 11940 9795 11996
rect 9795 11940 9799 11996
rect 9735 11936 9799 11940
rect 9815 11996 9879 12000
rect 9815 11940 9819 11996
rect 9819 11940 9875 11996
rect 9875 11940 9879 11996
rect 9815 11936 9879 11940
rect 9895 11996 9959 12000
rect 9895 11940 9899 11996
rect 9899 11940 9955 11996
rect 9955 11940 9959 11996
rect 9895 11936 9959 11940
rect 13357 11996 13421 12000
rect 13357 11940 13361 11996
rect 13361 11940 13417 11996
rect 13417 11940 13421 11996
rect 13357 11936 13421 11940
rect 13437 11996 13501 12000
rect 13437 11940 13441 11996
rect 13441 11940 13497 11996
rect 13497 11940 13501 11996
rect 13437 11936 13501 11940
rect 13517 11996 13581 12000
rect 13517 11940 13521 11996
rect 13521 11940 13577 11996
rect 13577 11940 13581 11996
rect 13517 11936 13581 11940
rect 13597 11996 13661 12000
rect 13597 11940 13601 11996
rect 13601 11940 13657 11996
rect 13657 11940 13661 11996
rect 13597 11936 13661 11940
rect 4102 11452 4166 11456
rect 4102 11396 4106 11452
rect 4106 11396 4162 11452
rect 4162 11396 4166 11452
rect 4102 11392 4166 11396
rect 4182 11452 4246 11456
rect 4182 11396 4186 11452
rect 4186 11396 4242 11452
rect 4242 11396 4246 11452
rect 4182 11392 4246 11396
rect 4262 11452 4326 11456
rect 4262 11396 4266 11452
rect 4266 11396 4322 11452
rect 4322 11396 4326 11452
rect 4262 11392 4326 11396
rect 4342 11452 4406 11456
rect 4342 11396 4346 11452
rect 4346 11396 4402 11452
rect 4402 11396 4406 11452
rect 4342 11392 4406 11396
rect 7804 11452 7868 11456
rect 7804 11396 7808 11452
rect 7808 11396 7864 11452
rect 7864 11396 7868 11452
rect 7804 11392 7868 11396
rect 7884 11452 7948 11456
rect 7884 11396 7888 11452
rect 7888 11396 7944 11452
rect 7944 11396 7948 11452
rect 7884 11392 7948 11396
rect 7964 11452 8028 11456
rect 7964 11396 7968 11452
rect 7968 11396 8024 11452
rect 8024 11396 8028 11452
rect 7964 11392 8028 11396
rect 8044 11452 8108 11456
rect 8044 11396 8048 11452
rect 8048 11396 8104 11452
rect 8104 11396 8108 11452
rect 8044 11392 8108 11396
rect 11506 11452 11570 11456
rect 11506 11396 11510 11452
rect 11510 11396 11566 11452
rect 11566 11396 11570 11452
rect 11506 11392 11570 11396
rect 11586 11452 11650 11456
rect 11586 11396 11590 11452
rect 11590 11396 11646 11452
rect 11646 11396 11650 11452
rect 11586 11392 11650 11396
rect 11666 11452 11730 11456
rect 11666 11396 11670 11452
rect 11670 11396 11726 11452
rect 11726 11396 11730 11452
rect 11666 11392 11730 11396
rect 11746 11452 11810 11456
rect 11746 11396 11750 11452
rect 11750 11396 11806 11452
rect 11806 11396 11810 11452
rect 11746 11392 11810 11396
rect 15208 11452 15272 11456
rect 15208 11396 15212 11452
rect 15212 11396 15268 11452
rect 15268 11396 15272 11452
rect 15208 11392 15272 11396
rect 15288 11452 15352 11456
rect 15288 11396 15292 11452
rect 15292 11396 15348 11452
rect 15348 11396 15352 11452
rect 15288 11392 15352 11396
rect 15368 11452 15432 11456
rect 15368 11396 15372 11452
rect 15372 11396 15428 11452
rect 15428 11396 15432 11452
rect 15368 11392 15432 11396
rect 15448 11452 15512 11456
rect 15448 11396 15452 11452
rect 15452 11396 15508 11452
rect 15508 11396 15512 11452
rect 15448 11392 15512 11396
rect 2251 10908 2315 10912
rect 2251 10852 2255 10908
rect 2255 10852 2311 10908
rect 2311 10852 2315 10908
rect 2251 10848 2315 10852
rect 2331 10908 2395 10912
rect 2331 10852 2335 10908
rect 2335 10852 2391 10908
rect 2391 10852 2395 10908
rect 2331 10848 2395 10852
rect 2411 10908 2475 10912
rect 2411 10852 2415 10908
rect 2415 10852 2471 10908
rect 2471 10852 2475 10908
rect 2411 10848 2475 10852
rect 2491 10908 2555 10912
rect 2491 10852 2495 10908
rect 2495 10852 2551 10908
rect 2551 10852 2555 10908
rect 2491 10848 2555 10852
rect 5953 10908 6017 10912
rect 5953 10852 5957 10908
rect 5957 10852 6013 10908
rect 6013 10852 6017 10908
rect 5953 10848 6017 10852
rect 6033 10908 6097 10912
rect 6033 10852 6037 10908
rect 6037 10852 6093 10908
rect 6093 10852 6097 10908
rect 6033 10848 6097 10852
rect 6113 10908 6177 10912
rect 6113 10852 6117 10908
rect 6117 10852 6173 10908
rect 6173 10852 6177 10908
rect 6113 10848 6177 10852
rect 6193 10908 6257 10912
rect 6193 10852 6197 10908
rect 6197 10852 6253 10908
rect 6253 10852 6257 10908
rect 6193 10848 6257 10852
rect 9655 10908 9719 10912
rect 9655 10852 9659 10908
rect 9659 10852 9715 10908
rect 9715 10852 9719 10908
rect 9655 10848 9719 10852
rect 9735 10908 9799 10912
rect 9735 10852 9739 10908
rect 9739 10852 9795 10908
rect 9795 10852 9799 10908
rect 9735 10848 9799 10852
rect 9815 10908 9879 10912
rect 9815 10852 9819 10908
rect 9819 10852 9875 10908
rect 9875 10852 9879 10908
rect 9815 10848 9879 10852
rect 9895 10908 9959 10912
rect 9895 10852 9899 10908
rect 9899 10852 9955 10908
rect 9955 10852 9959 10908
rect 9895 10848 9959 10852
rect 13357 10908 13421 10912
rect 13357 10852 13361 10908
rect 13361 10852 13417 10908
rect 13417 10852 13421 10908
rect 13357 10848 13421 10852
rect 13437 10908 13501 10912
rect 13437 10852 13441 10908
rect 13441 10852 13497 10908
rect 13497 10852 13501 10908
rect 13437 10848 13501 10852
rect 13517 10908 13581 10912
rect 13517 10852 13521 10908
rect 13521 10852 13577 10908
rect 13577 10852 13581 10908
rect 13517 10848 13581 10852
rect 13597 10908 13661 10912
rect 13597 10852 13601 10908
rect 13601 10852 13657 10908
rect 13657 10852 13661 10908
rect 13597 10848 13661 10852
rect 4102 10364 4166 10368
rect 4102 10308 4106 10364
rect 4106 10308 4162 10364
rect 4162 10308 4166 10364
rect 4102 10304 4166 10308
rect 4182 10364 4246 10368
rect 4182 10308 4186 10364
rect 4186 10308 4242 10364
rect 4242 10308 4246 10364
rect 4182 10304 4246 10308
rect 4262 10364 4326 10368
rect 4262 10308 4266 10364
rect 4266 10308 4322 10364
rect 4322 10308 4326 10364
rect 4262 10304 4326 10308
rect 4342 10364 4406 10368
rect 4342 10308 4346 10364
rect 4346 10308 4402 10364
rect 4402 10308 4406 10364
rect 4342 10304 4406 10308
rect 7804 10364 7868 10368
rect 7804 10308 7808 10364
rect 7808 10308 7864 10364
rect 7864 10308 7868 10364
rect 7804 10304 7868 10308
rect 7884 10364 7948 10368
rect 7884 10308 7888 10364
rect 7888 10308 7944 10364
rect 7944 10308 7948 10364
rect 7884 10304 7948 10308
rect 7964 10364 8028 10368
rect 7964 10308 7968 10364
rect 7968 10308 8024 10364
rect 8024 10308 8028 10364
rect 7964 10304 8028 10308
rect 8044 10364 8108 10368
rect 8044 10308 8048 10364
rect 8048 10308 8104 10364
rect 8104 10308 8108 10364
rect 8044 10304 8108 10308
rect 11506 10364 11570 10368
rect 11506 10308 11510 10364
rect 11510 10308 11566 10364
rect 11566 10308 11570 10364
rect 11506 10304 11570 10308
rect 11586 10364 11650 10368
rect 11586 10308 11590 10364
rect 11590 10308 11646 10364
rect 11646 10308 11650 10364
rect 11586 10304 11650 10308
rect 11666 10364 11730 10368
rect 11666 10308 11670 10364
rect 11670 10308 11726 10364
rect 11726 10308 11730 10364
rect 11666 10304 11730 10308
rect 11746 10364 11810 10368
rect 11746 10308 11750 10364
rect 11750 10308 11806 10364
rect 11806 10308 11810 10364
rect 11746 10304 11810 10308
rect 15208 10364 15272 10368
rect 15208 10308 15212 10364
rect 15212 10308 15268 10364
rect 15268 10308 15272 10364
rect 15208 10304 15272 10308
rect 15288 10364 15352 10368
rect 15288 10308 15292 10364
rect 15292 10308 15348 10364
rect 15348 10308 15352 10364
rect 15288 10304 15352 10308
rect 15368 10364 15432 10368
rect 15368 10308 15372 10364
rect 15372 10308 15428 10364
rect 15428 10308 15432 10364
rect 15368 10304 15432 10308
rect 15448 10364 15512 10368
rect 15448 10308 15452 10364
rect 15452 10308 15508 10364
rect 15508 10308 15512 10364
rect 15448 10304 15512 10308
rect 2251 9820 2315 9824
rect 2251 9764 2255 9820
rect 2255 9764 2311 9820
rect 2311 9764 2315 9820
rect 2251 9760 2315 9764
rect 2331 9820 2395 9824
rect 2331 9764 2335 9820
rect 2335 9764 2391 9820
rect 2391 9764 2395 9820
rect 2331 9760 2395 9764
rect 2411 9820 2475 9824
rect 2411 9764 2415 9820
rect 2415 9764 2471 9820
rect 2471 9764 2475 9820
rect 2411 9760 2475 9764
rect 2491 9820 2555 9824
rect 2491 9764 2495 9820
rect 2495 9764 2551 9820
rect 2551 9764 2555 9820
rect 2491 9760 2555 9764
rect 5953 9820 6017 9824
rect 5953 9764 5957 9820
rect 5957 9764 6013 9820
rect 6013 9764 6017 9820
rect 5953 9760 6017 9764
rect 6033 9820 6097 9824
rect 6033 9764 6037 9820
rect 6037 9764 6093 9820
rect 6093 9764 6097 9820
rect 6033 9760 6097 9764
rect 6113 9820 6177 9824
rect 6113 9764 6117 9820
rect 6117 9764 6173 9820
rect 6173 9764 6177 9820
rect 6113 9760 6177 9764
rect 6193 9820 6257 9824
rect 6193 9764 6197 9820
rect 6197 9764 6253 9820
rect 6253 9764 6257 9820
rect 6193 9760 6257 9764
rect 9655 9820 9719 9824
rect 9655 9764 9659 9820
rect 9659 9764 9715 9820
rect 9715 9764 9719 9820
rect 9655 9760 9719 9764
rect 9735 9820 9799 9824
rect 9735 9764 9739 9820
rect 9739 9764 9795 9820
rect 9795 9764 9799 9820
rect 9735 9760 9799 9764
rect 9815 9820 9879 9824
rect 9815 9764 9819 9820
rect 9819 9764 9875 9820
rect 9875 9764 9879 9820
rect 9815 9760 9879 9764
rect 9895 9820 9959 9824
rect 9895 9764 9899 9820
rect 9899 9764 9955 9820
rect 9955 9764 9959 9820
rect 9895 9760 9959 9764
rect 13357 9820 13421 9824
rect 13357 9764 13361 9820
rect 13361 9764 13417 9820
rect 13417 9764 13421 9820
rect 13357 9760 13421 9764
rect 13437 9820 13501 9824
rect 13437 9764 13441 9820
rect 13441 9764 13497 9820
rect 13497 9764 13501 9820
rect 13437 9760 13501 9764
rect 13517 9820 13581 9824
rect 13517 9764 13521 9820
rect 13521 9764 13577 9820
rect 13577 9764 13581 9820
rect 13517 9760 13581 9764
rect 13597 9820 13661 9824
rect 13597 9764 13601 9820
rect 13601 9764 13657 9820
rect 13657 9764 13661 9820
rect 13597 9760 13661 9764
rect 4102 9276 4166 9280
rect 4102 9220 4106 9276
rect 4106 9220 4162 9276
rect 4162 9220 4166 9276
rect 4102 9216 4166 9220
rect 4182 9276 4246 9280
rect 4182 9220 4186 9276
rect 4186 9220 4242 9276
rect 4242 9220 4246 9276
rect 4182 9216 4246 9220
rect 4262 9276 4326 9280
rect 4262 9220 4266 9276
rect 4266 9220 4322 9276
rect 4322 9220 4326 9276
rect 4262 9216 4326 9220
rect 4342 9276 4406 9280
rect 4342 9220 4346 9276
rect 4346 9220 4402 9276
rect 4402 9220 4406 9276
rect 4342 9216 4406 9220
rect 7804 9276 7868 9280
rect 7804 9220 7808 9276
rect 7808 9220 7864 9276
rect 7864 9220 7868 9276
rect 7804 9216 7868 9220
rect 7884 9276 7948 9280
rect 7884 9220 7888 9276
rect 7888 9220 7944 9276
rect 7944 9220 7948 9276
rect 7884 9216 7948 9220
rect 7964 9276 8028 9280
rect 7964 9220 7968 9276
rect 7968 9220 8024 9276
rect 8024 9220 8028 9276
rect 7964 9216 8028 9220
rect 8044 9276 8108 9280
rect 8044 9220 8048 9276
rect 8048 9220 8104 9276
rect 8104 9220 8108 9276
rect 8044 9216 8108 9220
rect 11506 9276 11570 9280
rect 11506 9220 11510 9276
rect 11510 9220 11566 9276
rect 11566 9220 11570 9276
rect 11506 9216 11570 9220
rect 11586 9276 11650 9280
rect 11586 9220 11590 9276
rect 11590 9220 11646 9276
rect 11646 9220 11650 9276
rect 11586 9216 11650 9220
rect 11666 9276 11730 9280
rect 11666 9220 11670 9276
rect 11670 9220 11726 9276
rect 11726 9220 11730 9276
rect 11666 9216 11730 9220
rect 11746 9276 11810 9280
rect 11746 9220 11750 9276
rect 11750 9220 11806 9276
rect 11806 9220 11810 9276
rect 11746 9216 11810 9220
rect 15208 9276 15272 9280
rect 15208 9220 15212 9276
rect 15212 9220 15268 9276
rect 15268 9220 15272 9276
rect 15208 9216 15272 9220
rect 15288 9276 15352 9280
rect 15288 9220 15292 9276
rect 15292 9220 15348 9276
rect 15348 9220 15352 9276
rect 15288 9216 15352 9220
rect 15368 9276 15432 9280
rect 15368 9220 15372 9276
rect 15372 9220 15428 9276
rect 15428 9220 15432 9276
rect 15368 9216 15432 9220
rect 15448 9276 15512 9280
rect 15448 9220 15452 9276
rect 15452 9220 15508 9276
rect 15508 9220 15512 9276
rect 15448 9216 15512 9220
rect 2251 8732 2315 8736
rect 2251 8676 2255 8732
rect 2255 8676 2311 8732
rect 2311 8676 2315 8732
rect 2251 8672 2315 8676
rect 2331 8732 2395 8736
rect 2331 8676 2335 8732
rect 2335 8676 2391 8732
rect 2391 8676 2395 8732
rect 2331 8672 2395 8676
rect 2411 8732 2475 8736
rect 2411 8676 2415 8732
rect 2415 8676 2471 8732
rect 2471 8676 2475 8732
rect 2411 8672 2475 8676
rect 2491 8732 2555 8736
rect 2491 8676 2495 8732
rect 2495 8676 2551 8732
rect 2551 8676 2555 8732
rect 2491 8672 2555 8676
rect 5953 8732 6017 8736
rect 5953 8676 5957 8732
rect 5957 8676 6013 8732
rect 6013 8676 6017 8732
rect 5953 8672 6017 8676
rect 6033 8732 6097 8736
rect 6033 8676 6037 8732
rect 6037 8676 6093 8732
rect 6093 8676 6097 8732
rect 6033 8672 6097 8676
rect 6113 8732 6177 8736
rect 6113 8676 6117 8732
rect 6117 8676 6173 8732
rect 6173 8676 6177 8732
rect 6113 8672 6177 8676
rect 6193 8732 6257 8736
rect 6193 8676 6197 8732
rect 6197 8676 6253 8732
rect 6253 8676 6257 8732
rect 6193 8672 6257 8676
rect 9655 8732 9719 8736
rect 9655 8676 9659 8732
rect 9659 8676 9715 8732
rect 9715 8676 9719 8732
rect 9655 8672 9719 8676
rect 9735 8732 9799 8736
rect 9735 8676 9739 8732
rect 9739 8676 9795 8732
rect 9795 8676 9799 8732
rect 9735 8672 9799 8676
rect 9815 8732 9879 8736
rect 9815 8676 9819 8732
rect 9819 8676 9875 8732
rect 9875 8676 9879 8732
rect 9815 8672 9879 8676
rect 9895 8732 9959 8736
rect 9895 8676 9899 8732
rect 9899 8676 9955 8732
rect 9955 8676 9959 8732
rect 9895 8672 9959 8676
rect 13357 8732 13421 8736
rect 13357 8676 13361 8732
rect 13361 8676 13417 8732
rect 13417 8676 13421 8732
rect 13357 8672 13421 8676
rect 13437 8732 13501 8736
rect 13437 8676 13441 8732
rect 13441 8676 13497 8732
rect 13497 8676 13501 8732
rect 13437 8672 13501 8676
rect 13517 8732 13581 8736
rect 13517 8676 13521 8732
rect 13521 8676 13577 8732
rect 13577 8676 13581 8732
rect 13517 8672 13581 8676
rect 13597 8732 13661 8736
rect 13597 8676 13601 8732
rect 13601 8676 13657 8732
rect 13657 8676 13661 8732
rect 13597 8672 13661 8676
rect 4102 8188 4166 8192
rect 4102 8132 4106 8188
rect 4106 8132 4162 8188
rect 4162 8132 4166 8188
rect 4102 8128 4166 8132
rect 4182 8188 4246 8192
rect 4182 8132 4186 8188
rect 4186 8132 4242 8188
rect 4242 8132 4246 8188
rect 4182 8128 4246 8132
rect 4262 8188 4326 8192
rect 4262 8132 4266 8188
rect 4266 8132 4322 8188
rect 4322 8132 4326 8188
rect 4262 8128 4326 8132
rect 4342 8188 4406 8192
rect 4342 8132 4346 8188
rect 4346 8132 4402 8188
rect 4402 8132 4406 8188
rect 4342 8128 4406 8132
rect 7804 8188 7868 8192
rect 7804 8132 7808 8188
rect 7808 8132 7864 8188
rect 7864 8132 7868 8188
rect 7804 8128 7868 8132
rect 7884 8188 7948 8192
rect 7884 8132 7888 8188
rect 7888 8132 7944 8188
rect 7944 8132 7948 8188
rect 7884 8128 7948 8132
rect 7964 8188 8028 8192
rect 7964 8132 7968 8188
rect 7968 8132 8024 8188
rect 8024 8132 8028 8188
rect 7964 8128 8028 8132
rect 8044 8188 8108 8192
rect 8044 8132 8048 8188
rect 8048 8132 8104 8188
rect 8104 8132 8108 8188
rect 8044 8128 8108 8132
rect 11506 8188 11570 8192
rect 11506 8132 11510 8188
rect 11510 8132 11566 8188
rect 11566 8132 11570 8188
rect 11506 8128 11570 8132
rect 11586 8188 11650 8192
rect 11586 8132 11590 8188
rect 11590 8132 11646 8188
rect 11646 8132 11650 8188
rect 11586 8128 11650 8132
rect 11666 8188 11730 8192
rect 11666 8132 11670 8188
rect 11670 8132 11726 8188
rect 11726 8132 11730 8188
rect 11666 8128 11730 8132
rect 11746 8188 11810 8192
rect 11746 8132 11750 8188
rect 11750 8132 11806 8188
rect 11806 8132 11810 8188
rect 11746 8128 11810 8132
rect 15208 8188 15272 8192
rect 15208 8132 15212 8188
rect 15212 8132 15268 8188
rect 15268 8132 15272 8188
rect 15208 8128 15272 8132
rect 15288 8188 15352 8192
rect 15288 8132 15292 8188
rect 15292 8132 15348 8188
rect 15348 8132 15352 8188
rect 15288 8128 15352 8132
rect 15368 8188 15432 8192
rect 15368 8132 15372 8188
rect 15372 8132 15428 8188
rect 15428 8132 15432 8188
rect 15368 8128 15432 8132
rect 15448 8188 15512 8192
rect 15448 8132 15452 8188
rect 15452 8132 15508 8188
rect 15508 8132 15512 8188
rect 15448 8128 15512 8132
rect 2251 7644 2315 7648
rect 2251 7588 2255 7644
rect 2255 7588 2311 7644
rect 2311 7588 2315 7644
rect 2251 7584 2315 7588
rect 2331 7644 2395 7648
rect 2331 7588 2335 7644
rect 2335 7588 2391 7644
rect 2391 7588 2395 7644
rect 2331 7584 2395 7588
rect 2411 7644 2475 7648
rect 2411 7588 2415 7644
rect 2415 7588 2471 7644
rect 2471 7588 2475 7644
rect 2411 7584 2475 7588
rect 2491 7644 2555 7648
rect 2491 7588 2495 7644
rect 2495 7588 2551 7644
rect 2551 7588 2555 7644
rect 2491 7584 2555 7588
rect 5953 7644 6017 7648
rect 5953 7588 5957 7644
rect 5957 7588 6013 7644
rect 6013 7588 6017 7644
rect 5953 7584 6017 7588
rect 6033 7644 6097 7648
rect 6033 7588 6037 7644
rect 6037 7588 6093 7644
rect 6093 7588 6097 7644
rect 6033 7584 6097 7588
rect 6113 7644 6177 7648
rect 6113 7588 6117 7644
rect 6117 7588 6173 7644
rect 6173 7588 6177 7644
rect 6113 7584 6177 7588
rect 6193 7644 6257 7648
rect 6193 7588 6197 7644
rect 6197 7588 6253 7644
rect 6253 7588 6257 7644
rect 6193 7584 6257 7588
rect 9655 7644 9719 7648
rect 9655 7588 9659 7644
rect 9659 7588 9715 7644
rect 9715 7588 9719 7644
rect 9655 7584 9719 7588
rect 9735 7644 9799 7648
rect 9735 7588 9739 7644
rect 9739 7588 9795 7644
rect 9795 7588 9799 7644
rect 9735 7584 9799 7588
rect 9815 7644 9879 7648
rect 9815 7588 9819 7644
rect 9819 7588 9875 7644
rect 9875 7588 9879 7644
rect 9815 7584 9879 7588
rect 9895 7644 9959 7648
rect 9895 7588 9899 7644
rect 9899 7588 9955 7644
rect 9955 7588 9959 7644
rect 9895 7584 9959 7588
rect 13357 7644 13421 7648
rect 13357 7588 13361 7644
rect 13361 7588 13417 7644
rect 13417 7588 13421 7644
rect 13357 7584 13421 7588
rect 13437 7644 13501 7648
rect 13437 7588 13441 7644
rect 13441 7588 13497 7644
rect 13497 7588 13501 7644
rect 13437 7584 13501 7588
rect 13517 7644 13581 7648
rect 13517 7588 13521 7644
rect 13521 7588 13577 7644
rect 13577 7588 13581 7644
rect 13517 7584 13581 7588
rect 13597 7644 13661 7648
rect 13597 7588 13601 7644
rect 13601 7588 13657 7644
rect 13657 7588 13661 7644
rect 13597 7584 13661 7588
rect 4102 7100 4166 7104
rect 4102 7044 4106 7100
rect 4106 7044 4162 7100
rect 4162 7044 4166 7100
rect 4102 7040 4166 7044
rect 4182 7100 4246 7104
rect 4182 7044 4186 7100
rect 4186 7044 4242 7100
rect 4242 7044 4246 7100
rect 4182 7040 4246 7044
rect 4262 7100 4326 7104
rect 4262 7044 4266 7100
rect 4266 7044 4322 7100
rect 4322 7044 4326 7100
rect 4262 7040 4326 7044
rect 4342 7100 4406 7104
rect 4342 7044 4346 7100
rect 4346 7044 4402 7100
rect 4402 7044 4406 7100
rect 4342 7040 4406 7044
rect 7804 7100 7868 7104
rect 7804 7044 7808 7100
rect 7808 7044 7864 7100
rect 7864 7044 7868 7100
rect 7804 7040 7868 7044
rect 7884 7100 7948 7104
rect 7884 7044 7888 7100
rect 7888 7044 7944 7100
rect 7944 7044 7948 7100
rect 7884 7040 7948 7044
rect 7964 7100 8028 7104
rect 7964 7044 7968 7100
rect 7968 7044 8024 7100
rect 8024 7044 8028 7100
rect 7964 7040 8028 7044
rect 8044 7100 8108 7104
rect 8044 7044 8048 7100
rect 8048 7044 8104 7100
rect 8104 7044 8108 7100
rect 8044 7040 8108 7044
rect 11506 7100 11570 7104
rect 11506 7044 11510 7100
rect 11510 7044 11566 7100
rect 11566 7044 11570 7100
rect 11506 7040 11570 7044
rect 11586 7100 11650 7104
rect 11586 7044 11590 7100
rect 11590 7044 11646 7100
rect 11646 7044 11650 7100
rect 11586 7040 11650 7044
rect 11666 7100 11730 7104
rect 11666 7044 11670 7100
rect 11670 7044 11726 7100
rect 11726 7044 11730 7100
rect 11666 7040 11730 7044
rect 11746 7100 11810 7104
rect 11746 7044 11750 7100
rect 11750 7044 11806 7100
rect 11806 7044 11810 7100
rect 11746 7040 11810 7044
rect 15208 7100 15272 7104
rect 15208 7044 15212 7100
rect 15212 7044 15268 7100
rect 15268 7044 15272 7100
rect 15208 7040 15272 7044
rect 15288 7100 15352 7104
rect 15288 7044 15292 7100
rect 15292 7044 15348 7100
rect 15348 7044 15352 7100
rect 15288 7040 15352 7044
rect 15368 7100 15432 7104
rect 15368 7044 15372 7100
rect 15372 7044 15428 7100
rect 15428 7044 15432 7100
rect 15368 7040 15432 7044
rect 15448 7100 15512 7104
rect 15448 7044 15452 7100
rect 15452 7044 15508 7100
rect 15508 7044 15512 7100
rect 15448 7040 15512 7044
rect 2251 6556 2315 6560
rect 2251 6500 2255 6556
rect 2255 6500 2311 6556
rect 2311 6500 2315 6556
rect 2251 6496 2315 6500
rect 2331 6556 2395 6560
rect 2331 6500 2335 6556
rect 2335 6500 2391 6556
rect 2391 6500 2395 6556
rect 2331 6496 2395 6500
rect 2411 6556 2475 6560
rect 2411 6500 2415 6556
rect 2415 6500 2471 6556
rect 2471 6500 2475 6556
rect 2411 6496 2475 6500
rect 2491 6556 2555 6560
rect 2491 6500 2495 6556
rect 2495 6500 2551 6556
rect 2551 6500 2555 6556
rect 2491 6496 2555 6500
rect 5953 6556 6017 6560
rect 5953 6500 5957 6556
rect 5957 6500 6013 6556
rect 6013 6500 6017 6556
rect 5953 6496 6017 6500
rect 6033 6556 6097 6560
rect 6033 6500 6037 6556
rect 6037 6500 6093 6556
rect 6093 6500 6097 6556
rect 6033 6496 6097 6500
rect 6113 6556 6177 6560
rect 6113 6500 6117 6556
rect 6117 6500 6173 6556
rect 6173 6500 6177 6556
rect 6113 6496 6177 6500
rect 6193 6556 6257 6560
rect 6193 6500 6197 6556
rect 6197 6500 6253 6556
rect 6253 6500 6257 6556
rect 6193 6496 6257 6500
rect 9655 6556 9719 6560
rect 9655 6500 9659 6556
rect 9659 6500 9715 6556
rect 9715 6500 9719 6556
rect 9655 6496 9719 6500
rect 9735 6556 9799 6560
rect 9735 6500 9739 6556
rect 9739 6500 9795 6556
rect 9795 6500 9799 6556
rect 9735 6496 9799 6500
rect 9815 6556 9879 6560
rect 9815 6500 9819 6556
rect 9819 6500 9875 6556
rect 9875 6500 9879 6556
rect 9815 6496 9879 6500
rect 9895 6556 9959 6560
rect 9895 6500 9899 6556
rect 9899 6500 9955 6556
rect 9955 6500 9959 6556
rect 9895 6496 9959 6500
rect 13357 6556 13421 6560
rect 13357 6500 13361 6556
rect 13361 6500 13417 6556
rect 13417 6500 13421 6556
rect 13357 6496 13421 6500
rect 13437 6556 13501 6560
rect 13437 6500 13441 6556
rect 13441 6500 13497 6556
rect 13497 6500 13501 6556
rect 13437 6496 13501 6500
rect 13517 6556 13581 6560
rect 13517 6500 13521 6556
rect 13521 6500 13577 6556
rect 13577 6500 13581 6556
rect 13517 6496 13581 6500
rect 13597 6556 13661 6560
rect 13597 6500 13601 6556
rect 13601 6500 13657 6556
rect 13657 6500 13661 6556
rect 13597 6496 13661 6500
rect 4102 6012 4166 6016
rect 4102 5956 4106 6012
rect 4106 5956 4162 6012
rect 4162 5956 4166 6012
rect 4102 5952 4166 5956
rect 4182 6012 4246 6016
rect 4182 5956 4186 6012
rect 4186 5956 4242 6012
rect 4242 5956 4246 6012
rect 4182 5952 4246 5956
rect 4262 6012 4326 6016
rect 4262 5956 4266 6012
rect 4266 5956 4322 6012
rect 4322 5956 4326 6012
rect 4262 5952 4326 5956
rect 4342 6012 4406 6016
rect 4342 5956 4346 6012
rect 4346 5956 4402 6012
rect 4402 5956 4406 6012
rect 4342 5952 4406 5956
rect 7804 6012 7868 6016
rect 7804 5956 7808 6012
rect 7808 5956 7864 6012
rect 7864 5956 7868 6012
rect 7804 5952 7868 5956
rect 7884 6012 7948 6016
rect 7884 5956 7888 6012
rect 7888 5956 7944 6012
rect 7944 5956 7948 6012
rect 7884 5952 7948 5956
rect 7964 6012 8028 6016
rect 7964 5956 7968 6012
rect 7968 5956 8024 6012
rect 8024 5956 8028 6012
rect 7964 5952 8028 5956
rect 8044 6012 8108 6016
rect 8044 5956 8048 6012
rect 8048 5956 8104 6012
rect 8104 5956 8108 6012
rect 8044 5952 8108 5956
rect 11506 6012 11570 6016
rect 11506 5956 11510 6012
rect 11510 5956 11566 6012
rect 11566 5956 11570 6012
rect 11506 5952 11570 5956
rect 11586 6012 11650 6016
rect 11586 5956 11590 6012
rect 11590 5956 11646 6012
rect 11646 5956 11650 6012
rect 11586 5952 11650 5956
rect 11666 6012 11730 6016
rect 11666 5956 11670 6012
rect 11670 5956 11726 6012
rect 11726 5956 11730 6012
rect 11666 5952 11730 5956
rect 11746 6012 11810 6016
rect 11746 5956 11750 6012
rect 11750 5956 11806 6012
rect 11806 5956 11810 6012
rect 11746 5952 11810 5956
rect 15208 6012 15272 6016
rect 15208 5956 15212 6012
rect 15212 5956 15268 6012
rect 15268 5956 15272 6012
rect 15208 5952 15272 5956
rect 15288 6012 15352 6016
rect 15288 5956 15292 6012
rect 15292 5956 15348 6012
rect 15348 5956 15352 6012
rect 15288 5952 15352 5956
rect 15368 6012 15432 6016
rect 15368 5956 15372 6012
rect 15372 5956 15428 6012
rect 15428 5956 15432 6012
rect 15368 5952 15432 5956
rect 15448 6012 15512 6016
rect 15448 5956 15452 6012
rect 15452 5956 15508 6012
rect 15508 5956 15512 6012
rect 15448 5952 15512 5956
rect 2251 5468 2315 5472
rect 2251 5412 2255 5468
rect 2255 5412 2311 5468
rect 2311 5412 2315 5468
rect 2251 5408 2315 5412
rect 2331 5468 2395 5472
rect 2331 5412 2335 5468
rect 2335 5412 2391 5468
rect 2391 5412 2395 5468
rect 2331 5408 2395 5412
rect 2411 5468 2475 5472
rect 2411 5412 2415 5468
rect 2415 5412 2471 5468
rect 2471 5412 2475 5468
rect 2411 5408 2475 5412
rect 2491 5468 2555 5472
rect 2491 5412 2495 5468
rect 2495 5412 2551 5468
rect 2551 5412 2555 5468
rect 2491 5408 2555 5412
rect 5953 5468 6017 5472
rect 5953 5412 5957 5468
rect 5957 5412 6013 5468
rect 6013 5412 6017 5468
rect 5953 5408 6017 5412
rect 6033 5468 6097 5472
rect 6033 5412 6037 5468
rect 6037 5412 6093 5468
rect 6093 5412 6097 5468
rect 6033 5408 6097 5412
rect 6113 5468 6177 5472
rect 6113 5412 6117 5468
rect 6117 5412 6173 5468
rect 6173 5412 6177 5468
rect 6113 5408 6177 5412
rect 6193 5468 6257 5472
rect 6193 5412 6197 5468
rect 6197 5412 6253 5468
rect 6253 5412 6257 5468
rect 6193 5408 6257 5412
rect 9655 5468 9719 5472
rect 9655 5412 9659 5468
rect 9659 5412 9715 5468
rect 9715 5412 9719 5468
rect 9655 5408 9719 5412
rect 9735 5468 9799 5472
rect 9735 5412 9739 5468
rect 9739 5412 9795 5468
rect 9795 5412 9799 5468
rect 9735 5408 9799 5412
rect 9815 5468 9879 5472
rect 9815 5412 9819 5468
rect 9819 5412 9875 5468
rect 9875 5412 9879 5468
rect 9815 5408 9879 5412
rect 9895 5468 9959 5472
rect 9895 5412 9899 5468
rect 9899 5412 9955 5468
rect 9955 5412 9959 5468
rect 9895 5408 9959 5412
rect 13357 5468 13421 5472
rect 13357 5412 13361 5468
rect 13361 5412 13417 5468
rect 13417 5412 13421 5468
rect 13357 5408 13421 5412
rect 13437 5468 13501 5472
rect 13437 5412 13441 5468
rect 13441 5412 13497 5468
rect 13497 5412 13501 5468
rect 13437 5408 13501 5412
rect 13517 5468 13581 5472
rect 13517 5412 13521 5468
rect 13521 5412 13577 5468
rect 13577 5412 13581 5468
rect 13517 5408 13581 5412
rect 13597 5468 13661 5472
rect 13597 5412 13601 5468
rect 13601 5412 13657 5468
rect 13657 5412 13661 5468
rect 13597 5408 13661 5412
rect 4102 4924 4166 4928
rect 4102 4868 4106 4924
rect 4106 4868 4162 4924
rect 4162 4868 4166 4924
rect 4102 4864 4166 4868
rect 4182 4924 4246 4928
rect 4182 4868 4186 4924
rect 4186 4868 4242 4924
rect 4242 4868 4246 4924
rect 4182 4864 4246 4868
rect 4262 4924 4326 4928
rect 4262 4868 4266 4924
rect 4266 4868 4322 4924
rect 4322 4868 4326 4924
rect 4262 4864 4326 4868
rect 4342 4924 4406 4928
rect 4342 4868 4346 4924
rect 4346 4868 4402 4924
rect 4402 4868 4406 4924
rect 4342 4864 4406 4868
rect 7804 4924 7868 4928
rect 7804 4868 7808 4924
rect 7808 4868 7864 4924
rect 7864 4868 7868 4924
rect 7804 4864 7868 4868
rect 7884 4924 7948 4928
rect 7884 4868 7888 4924
rect 7888 4868 7944 4924
rect 7944 4868 7948 4924
rect 7884 4864 7948 4868
rect 7964 4924 8028 4928
rect 7964 4868 7968 4924
rect 7968 4868 8024 4924
rect 8024 4868 8028 4924
rect 7964 4864 8028 4868
rect 8044 4924 8108 4928
rect 8044 4868 8048 4924
rect 8048 4868 8104 4924
rect 8104 4868 8108 4924
rect 8044 4864 8108 4868
rect 11506 4924 11570 4928
rect 11506 4868 11510 4924
rect 11510 4868 11566 4924
rect 11566 4868 11570 4924
rect 11506 4864 11570 4868
rect 11586 4924 11650 4928
rect 11586 4868 11590 4924
rect 11590 4868 11646 4924
rect 11646 4868 11650 4924
rect 11586 4864 11650 4868
rect 11666 4924 11730 4928
rect 11666 4868 11670 4924
rect 11670 4868 11726 4924
rect 11726 4868 11730 4924
rect 11666 4864 11730 4868
rect 11746 4924 11810 4928
rect 11746 4868 11750 4924
rect 11750 4868 11806 4924
rect 11806 4868 11810 4924
rect 11746 4864 11810 4868
rect 15208 4924 15272 4928
rect 15208 4868 15212 4924
rect 15212 4868 15268 4924
rect 15268 4868 15272 4924
rect 15208 4864 15272 4868
rect 15288 4924 15352 4928
rect 15288 4868 15292 4924
rect 15292 4868 15348 4924
rect 15348 4868 15352 4924
rect 15288 4864 15352 4868
rect 15368 4924 15432 4928
rect 15368 4868 15372 4924
rect 15372 4868 15428 4924
rect 15428 4868 15432 4924
rect 15368 4864 15432 4868
rect 15448 4924 15512 4928
rect 15448 4868 15452 4924
rect 15452 4868 15508 4924
rect 15508 4868 15512 4924
rect 15448 4864 15512 4868
rect 2251 4380 2315 4384
rect 2251 4324 2255 4380
rect 2255 4324 2311 4380
rect 2311 4324 2315 4380
rect 2251 4320 2315 4324
rect 2331 4380 2395 4384
rect 2331 4324 2335 4380
rect 2335 4324 2391 4380
rect 2391 4324 2395 4380
rect 2331 4320 2395 4324
rect 2411 4380 2475 4384
rect 2411 4324 2415 4380
rect 2415 4324 2471 4380
rect 2471 4324 2475 4380
rect 2411 4320 2475 4324
rect 2491 4380 2555 4384
rect 2491 4324 2495 4380
rect 2495 4324 2551 4380
rect 2551 4324 2555 4380
rect 2491 4320 2555 4324
rect 5953 4380 6017 4384
rect 5953 4324 5957 4380
rect 5957 4324 6013 4380
rect 6013 4324 6017 4380
rect 5953 4320 6017 4324
rect 6033 4380 6097 4384
rect 6033 4324 6037 4380
rect 6037 4324 6093 4380
rect 6093 4324 6097 4380
rect 6033 4320 6097 4324
rect 6113 4380 6177 4384
rect 6113 4324 6117 4380
rect 6117 4324 6173 4380
rect 6173 4324 6177 4380
rect 6113 4320 6177 4324
rect 6193 4380 6257 4384
rect 6193 4324 6197 4380
rect 6197 4324 6253 4380
rect 6253 4324 6257 4380
rect 6193 4320 6257 4324
rect 9655 4380 9719 4384
rect 9655 4324 9659 4380
rect 9659 4324 9715 4380
rect 9715 4324 9719 4380
rect 9655 4320 9719 4324
rect 9735 4380 9799 4384
rect 9735 4324 9739 4380
rect 9739 4324 9795 4380
rect 9795 4324 9799 4380
rect 9735 4320 9799 4324
rect 9815 4380 9879 4384
rect 9815 4324 9819 4380
rect 9819 4324 9875 4380
rect 9875 4324 9879 4380
rect 9815 4320 9879 4324
rect 9895 4380 9959 4384
rect 9895 4324 9899 4380
rect 9899 4324 9955 4380
rect 9955 4324 9959 4380
rect 9895 4320 9959 4324
rect 13357 4380 13421 4384
rect 13357 4324 13361 4380
rect 13361 4324 13417 4380
rect 13417 4324 13421 4380
rect 13357 4320 13421 4324
rect 13437 4380 13501 4384
rect 13437 4324 13441 4380
rect 13441 4324 13497 4380
rect 13497 4324 13501 4380
rect 13437 4320 13501 4324
rect 13517 4380 13581 4384
rect 13517 4324 13521 4380
rect 13521 4324 13577 4380
rect 13577 4324 13581 4380
rect 13517 4320 13581 4324
rect 13597 4380 13661 4384
rect 13597 4324 13601 4380
rect 13601 4324 13657 4380
rect 13657 4324 13661 4380
rect 13597 4320 13661 4324
rect 4102 3836 4166 3840
rect 4102 3780 4106 3836
rect 4106 3780 4162 3836
rect 4162 3780 4166 3836
rect 4102 3776 4166 3780
rect 4182 3836 4246 3840
rect 4182 3780 4186 3836
rect 4186 3780 4242 3836
rect 4242 3780 4246 3836
rect 4182 3776 4246 3780
rect 4262 3836 4326 3840
rect 4262 3780 4266 3836
rect 4266 3780 4322 3836
rect 4322 3780 4326 3836
rect 4262 3776 4326 3780
rect 4342 3836 4406 3840
rect 4342 3780 4346 3836
rect 4346 3780 4402 3836
rect 4402 3780 4406 3836
rect 4342 3776 4406 3780
rect 7804 3836 7868 3840
rect 7804 3780 7808 3836
rect 7808 3780 7864 3836
rect 7864 3780 7868 3836
rect 7804 3776 7868 3780
rect 7884 3836 7948 3840
rect 7884 3780 7888 3836
rect 7888 3780 7944 3836
rect 7944 3780 7948 3836
rect 7884 3776 7948 3780
rect 7964 3836 8028 3840
rect 7964 3780 7968 3836
rect 7968 3780 8024 3836
rect 8024 3780 8028 3836
rect 7964 3776 8028 3780
rect 8044 3836 8108 3840
rect 8044 3780 8048 3836
rect 8048 3780 8104 3836
rect 8104 3780 8108 3836
rect 8044 3776 8108 3780
rect 11506 3836 11570 3840
rect 11506 3780 11510 3836
rect 11510 3780 11566 3836
rect 11566 3780 11570 3836
rect 11506 3776 11570 3780
rect 11586 3836 11650 3840
rect 11586 3780 11590 3836
rect 11590 3780 11646 3836
rect 11646 3780 11650 3836
rect 11586 3776 11650 3780
rect 11666 3836 11730 3840
rect 11666 3780 11670 3836
rect 11670 3780 11726 3836
rect 11726 3780 11730 3836
rect 11666 3776 11730 3780
rect 11746 3836 11810 3840
rect 11746 3780 11750 3836
rect 11750 3780 11806 3836
rect 11806 3780 11810 3836
rect 11746 3776 11810 3780
rect 15208 3836 15272 3840
rect 15208 3780 15212 3836
rect 15212 3780 15268 3836
rect 15268 3780 15272 3836
rect 15208 3776 15272 3780
rect 15288 3836 15352 3840
rect 15288 3780 15292 3836
rect 15292 3780 15348 3836
rect 15348 3780 15352 3836
rect 15288 3776 15352 3780
rect 15368 3836 15432 3840
rect 15368 3780 15372 3836
rect 15372 3780 15428 3836
rect 15428 3780 15432 3836
rect 15368 3776 15432 3780
rect 15448 3836 15512 3840
rect 15448 3780 15452 3836
rect 15452 3780 15508 3836
rect 15508 3780 15512 3836
rect 15448 3776 15512 3780
rect 2251 3292 2315 3296
rect 2251 3236 2255 3292
rect 2255 3236 2311 3292
rect 2311 3236 2315 3292
rect 2251 3232 2315 3236
rect 2331 3292 2395 3296
rect 2331 3236 2335 3292
rect 2335 3236 2391 3292
rect 2391 3236 2395 3292
rect 2331 3232 2395 3236
rect 2411 3292 2475 3296
rect 2411 3236 2415 3292
rect 2415 3236 2471 3292
rect 2471 3236 2475 3292
rect 2411 3232 2475 3236
rect 2491 3292 2555 3296
rect 2491 3236 2495 3292
rect 2495 3236 2551 3292
rect 2551 3236 2555 3292
rect 2491 3232 2555 3236
rect 5953 3292 6017 3296
rect 5953 3236 5957 3292
rect 5957 3236 6013 3292
rect 6013 3236 6017 3292
rect 5953 3232 6017 3236
rect 6033 3292 6097 3296
rect 6033 3236 6037 3292
rect 6037 3236 6093 3292
rect 6093 3236 6097 3292
rect 6033 3232 6097 3236
rect 6113 3292 6177 3296
rect 6113 3236 6117 3292
rect 6117 3236 6173 3292
rect 6173 3236 6177 3292
rect 6113 3232 6177 3236
rect 6193 3292 6257 3296
rect 6193 3236 6197 3292
rect 6197 3236 6253 3292
rect 6253 3236 6257 3292
rect 6193 3232 6257 3236
rect 9655 3292 9719 3296
rect 9655 3236 9659 3292
rect 9659 3236 9715 3292
rect 9715 3236 9719 3292
rect 9655 3232 9719 3236
rect 9735 3292 9799 3296
rect 9735 3236 9739 3292
rect 9739 3236 9795 3292
rect 9795 3236 9799 3292
rect 9735 3232 9799 3236
rect 9815 3292 9879 3296
rect 9815 3236 9819 3292
rect 9819 3236 9875 3292
rect 9875 3236 9879 3292
rect 9815 3232 9879 3236
rect 9895 3292 9959 3296
rect 9895 3236 9899 3292
rect 9899 3236 9955 3292
rect 9955 3236 9959 3292
rect 9895 3232 9959 3236
rect 13357 3292 13421 3296
rect 13357 3236 13361 3292
rect 13361 3236 13417 3292
rect 13417 3236 13421 3292
rect 13357 3232 13421 3236
rect 13437 3292 13501 3296
rect 13437 3236 13441 3292
rect 13441 3236 13497 3292
rect 13497 3236 13501 3292
rect 13437 3232 13501 3236
rect 13517 3292 13581 3296
rect 13517 3236 13521 3292
rect 13521 3236 13577 3292
rect 13577 3236 13581 3292
rect 13517 3232 13581 3236
rect 13597 3292 13661 3296
rect 13597 3236 13601 3292
rect 13601 3236 13657 3292
rect 13657 3236 13661 3292
rect 13597 3232 13661 3236
rect 4102 2748 4166 2752
rect 4102 2692 4106 2748
rect 4106 2692 4162 2748
rect 4162 2692 4166 2748
rect 4102 2688 4166 2692
rect 4182 2748 4246 2752
rect 4182 2692 4186 2748
rect 4186 2692 4242 2748
rect 4242 2692 4246 2748
rect 4182 2688 4246 2692
rect 4262 2748 4326 2752
rect 4262 2692 4266 2748
rect 4266 2692 4322 2748
rect 4322 2692 4326 2748
rect 4262 2688 4326 2692
rect 4342 2748 4406 2752
rect 4342 2692 4346 2748
rect 4346 2692 4402 2748
rect 4402 2692 4406 2748
rect 4342 2688 4406 2692
rect 7804 2748 7868 2752
rect 7804 2692 7808 2748
rect 7808 2692 7864 2748
rect 7864 2692 7868 2748
rect 7804 2688 7868 2692
rect 7884 2748 7948 2752
rect 7884 2692 7888 2748
rect 7888 2692 7944 2748
rect 7944 2692 7948 2748
rect 7884 2688 7948 2692
rect 7964 2748 8028 2752
rect 7964 2692 7968 2748
rect 7968 2692 8024 2748
rect 8024 2692 8028 2748
rect 7964 2688 8028 2692
rect 8044 2748 8108 2752
rect 8044 2692 8048 2748
rect 8048 2692 8104 2748
rect 8104 2692 8108 2748
rect 8044 2688 8108 2692
rect 11506 2748 11570 2752
rect 11506 2692 11510 2748
rect 11510 2692 11566 2748
rect 11566 2692 11570 2748
rect 11506 2688 11570 2692
rect 11586 2748 11650 2752
rect 11586 2692 11590 2748
rect 11590 2692 11646 2748
rect 11646 2692 11650 2748
rect 11586 2688 11650 2692
rect 11666 2748 11730 2752
rect 11666 2692 11670 2748
rect 11670 2692 11726 2748
rect 11726 2692 11730 2748
rect 11666 2688 11730 2692
rect 11746 2748 11810 2752
rect 11746 2692 11750 2748
rect 11750 2692 11806 2748
rect 11806 2692 11810 2748
rect 11746 2688 11810 2692
rect 15208 2748 15272 2752
rect 15208 2692 15212 2748
rect 15212 2692 15268 2748
rect 15268 2692 15272 2748
rect 15208 2688 15272 2692
rect 15288 2748 15352 2752
rect 15288 2692 15292 2748
rect 15292 2692 15348 2748
rect 15348 2692 15352 2748
rect 15288 2688 15352 2692
rect 15368 2748 15432 2752
rect 15368 2692 15372 2748
rect 15372 2692 15428 2748
rect 15428 2692 15432 2748
rect 15368 2688 15432 2692
rect 15448 2748 15512 2752
rect 15448 2692 15452 2748
rect 15452 2692 15508 2748
rect 15508 2692 15512 2748
rect 15448 2688 15512 2692
rect 2251 2204 2315 2208
rect 2251 2148 2255 2204
rect 2255 2148 2311 2204
rect 2311 2148 2315 2204
rect 2251 2144 2315 2148
rect 2331 2204 2395 2208
rect 2331 2148 2335 2204
rect 2335 2148 2391 2204
rect 2391 2148 2395 2204
rect 2331 2144 2395 2148
rect 2411 2204 2475 2208
rect 2411 2148 2415 2204
rect 2415 2148 2471 2204
rect 2471 2148 2475 2204
rect 2411 2144 2475 2148
rect 2491 2204 2555 2208
rect 2491 2148 2495 2204
rect 2495 2148 2551 2204
rect 2551 2148 2555 2204
rect 2491 2144 2555 2148
rect 5953 2204 6017 2208
rect 5953 2148 5957 2204
rect 5957 2148 6013 2204
rect 6013 2148 6017 2204
rect 5953 2144 6017 2148
rect 6033 2204 6097 2208
rect 6033 2148 6037 2204
rect 6037 2148 6093 2204
rect 6093 2148 6097 2204
rect 6033 2144 6097 2148
rect 6113 2204 6177 2208
rect 6113 2148 6117 2204
rect 6117 2148 6173 2204
rect 6173 2148 6177 2204
rect 6113 2144 6177 2148
rect 6193 2204 6257 2208
rect 6193 2148 6197 2204
rect 6197 2148 6253 2204
rect 6253 2148 6257 2204
rect 6193 2144 6257 2148
rect 9655 2204 9719 2208
rect 9655 2148 9659 2204
rect 9659 2148 9715 2204
rect 9715 2148 9719 2204
rect 9655 2144 9719 2148
rect 9735 2204 9799 2208
rect 9735 2148 9739 2204
rect 9739 2148 9795 2204
rect 9795 2148 9799 2204
rect 9735 2144 9799 2148
rect 9815 2204 9879 2208
rect 9815 2148 9819 2204
rect 9819 2148 9875 2204
rect 9875 2148 9879 2204
rect 9815 2144 9879 2148
rect 9895 2204 9959 2208
rect 9895 2148 9899 2204
rect 9899 2148 9955 2204
rect 9955 2148 9959 2204
rect 9895 2144 9959 2148
rect 13357 2204 13421 2208
rect 13357 2148 13361 2204
rect 13361 2148 13417 2204
rect 13417 2148 13421 2204
rect 13357 2144 13421 2148
rect 13437 2204 13501 2208
rect 13437 2148 13441 2204
rect 13441 2148 13497 2204
rect 13497 2148 13501 2204
rect 13437 2144 13501 2148
rect 13517 2204 13581 2208
rect 13517 2148 13521 2204
rect 13521 2148 13577 2204
rect 13577 2148 13581 2204
rect 13517 2144 13581 2148
rect 13597 2204 13661 2208
rect 13597 2148 13601 2204
rect 13601 2148 13657 2204
rect 13657 2148 13661 2204
rect 13597 2144 13661 2148
rect 4102 1660 4166 1664
rect 4102 1604 4106 1660
rect 4106 1604 4162 1660
rect 4162 1604 4166 1660
rect 4102 1600 4166 1604
rect 4182 1660 4246 1664
rect 4182 1604 4186 1660
rect 4186 1604 4242 1660
rect 4242 1604 4246 1660
rect 4182 1600 4246 1604
rect 4262 1660 4326 1664
rect 4262 1604 4266 1660
rect 4266 1604 4322 1660
rect 4322 1604 4326 1660
rect 4262 1600 4326 1604
rect 4342 1660 4406 1664
rect 4342 1604 4346 1660
rect 4346 1604 4402 1660
rect 4402 1604 4406 1660
rect 4342 1600 4406 1604
rect 7804 1660 7868 1664
rect 7804 1604 7808 1660
rect 7808 1604 7864 1660
rect 7864 1604 7868 1660
rect 7804 1600 7868 1604
rect 7884 1660 7948 1664
rect 7884 1604 7888 1660
rect 7888 1604 7944 1660
rect 7944 1604 7948 1660
rect 7884 1600 7948 1604
rect 7964 1660 8028 1664
rect 7964 1604 7968 1660
rect 7968 1604 8024 1660
rect 8024 1604 8028 1660
rect 7964 1600 8028 1604
rect 8044 1660 8108 1664
rect 8044 1604 8048 1660
rect 8048 1604 8104 1660
rect 8104 1604 8108 1660
rect 8044 1600 8108 1604
rect 11506 1660 11570 1664
rect 11506 1604 11510 1660
rect 11510 1604 11566 1660
rect 11566 1604 11570 1660
rect 11506 1600 11570 1604
rect 11586 1660 11650 1664
rect 11586 1604 11590 1660
rect 11590 1604 11646 1660
rect 11646 1604 11650 1660
rect 11586 1600 11650 1604
rect 11666 1660 11730 1664
rect 11666 1604 11670 1660
rect 11670 1604 11726 1660
rect 11726 1604 11730 1660
rect 11666 1600 11730 1604
rect 11746 1660 11810 1664
rect 11746 1604 11750 1660
rect 11750 1604 11806 1660
rect 11806 1604 11810 1660
rect 11746 1600 11810 1604
rect 15208 1660 15272 1664
rect 15208 1604 15212 1660
rect 15212 1604 15268 1660
rect 15268 1604 15272 1660
rect 15208 1600 15272 1604
rect 15288 1660 15352 1664
rect 15288 1604 15292 1660
rect 15292 1604 15348 1660
rect 15348 1604 15352 1660
rect 15288 1600 15352 1604
rect 15368 1660 15432 1664
rect 15368 1604 15372 1660
rect 15372 1604 15428 1660
rect 15428 1604 15432 1660
rect 15368 1600 15432 1604
rect 15448 1660 15512 1664
rect 15448 1604 15452 1660
rect 15452 1604 15508 1660
rect 15508 1604 15512 1660
rect 15448 1600 15512 1604
rect 2251 1116 2315 1120
rect 2251 1060 2255 1116
rect 2255 1060 2311 1116
rect 2311 1060 2315 1116
rect 2251 1056 2315 1060
rect 2331 1116 2395 1120
rect 2331 1060 2335 1116
rect 2335 1060 2391 1116
rect 2391 1060 2395 1116
rect 2331 1056 2395 1060
rect 2411 1116 2475 1120
rect 2411 1060 2415 1116
rect 2415 1060 2471 1116
rect 2471 1060 2475 1116
rect 2411 1056 2475 1060
rect 2491 1116 2555 1120
rect 2491 1060 2495 1116
rect 2495 1060 2551 1116
rect 2551 1060 2555 1116
rect 2491 1056 2555 1060
rect 5953 1116 6017 1120
rect 5953 1060 5957 1116
rect 5957 1060 6013 1116
rect 6013 1060 6017 1116
rect 5953 1056 6017 1060
rect 6033 1116 6097 1120
rect 6033 1060 6037 1116
rect 6037 1060 6093 1116
rect 6093 1060 6097 1116
rect 6033 1056 6097 1060
rect 6113 1116 6177 1120
rect 6113 1060 6117 1116
rect 6117 1060 6173 1116
rect 6173 1060 6177 1116
rect 6113 1056 6177 1060
rect 6193 1116 6257 1120
rect 6193 1060 6197 1116
rect 6197 1060 6253 1116
rect 6253 1060 6257 1116
rect 6193 1056 6257 1060
rect 9655 1116 9719 1120
rect 9655 1060 9659 1116
rect 9659 1060 9715 1116
rect 9715 1060 9719 1116
rect 9655 1056 9719 1060
rect 9735 1116 9799 1120
rect 9735 1060 9739 1116
rect 9739 1060 9795 1116
rect 9795 1060 9799 1116
rect 9735 1056 9799 1060
rect 9815 1116 9879 1120
rect 9815 1060 9819 1116
rect 9819 1060 9875 1116
rect 9875 1060 9879 1116
rect 9815 1056 9879 1060
rect 9895 1116 9959 1120
rect 9895 1060 9899 1116
rect 9899 1060 9955 1116
rect 9955 1060 9959 1116
rect 9895 1056 9959 1060
rect 13357 1116 13421 1120
rect 13357 1060 13361 1116
rect 13361 1060 13417 1116
rect 13417 1060 13421 1116
rect 13357 1056 13421 1060
rect 13437 1116 13501 1120
rect 13437 1060 13441 1116
rect 13441 1060 13497 1116
rect 13497 1060 13501 1116
rect 13437 1056 13501 1060
rect 13517 1116 13581 1120
rect 13517 1060 13521 1116
rect 13521 1060 13577 1116
rect 13577 1060 13581 1116
rect 13517 1056 13581 1060
rect 13597 1116 13661 1120
rect 13597 1060 13601 1116
rect 13601 1060 13657 1116
rect 13657 1060 13661 1116
rect 13597 1056 13661 1060
rect 4102 572 4166 576
rect 4102 516 4106 572
rect 4106 516 4162 572
rect 4162 516 4166 572
rect 4102 512 4166 516
rect 4182 572 4246 576
rect 4182 516 4186 572
rect 4186 516 4242 572
rect 4242 516 4246 572
rect 4182 512 4246 516
rect 4262 572 4326 576
rect 4262 516 4266 572
rect 4266 516 4322 572
rect 4322 516 4326 572
rect 4262 512 4326 516
rect 4342 572 4406 576
rect 4342 516 4346 572
rect 4346 516 4402 572
rect 4402 516 4406 572
rect 4342 512 4406 516
rect 7804 572 7868 576
rect 7804 516 7808 572
rect 7808 516 7864 572
rect 7864 516 7868 572
rect 7804 512 7868 516
rect 7884 572 7948 576
rect 7884 516 7888 572
rect 7888 516 7944 572
rect 7944 516 7948 572
rect 7884 512 7948 516
rect 7964 572 8028 576
rect 7964 516 7968 572
rect 7968 516 8024 572
rect 8024 516 8028 572
rect 7964 512 8028 516
rect 8044 572 8108 576
rect 8044 516 8048 572
rect 8048 516 8104 572
rect 8104 516 8108 572
rect 8044 512 8108 516
rect 11506 572 11570 576
rect 11506 516 11510 572
rect 11510 516 11566 572
rect 11566 516 11570 572
rect 11506 512 11570 516
rect 11586 572 11650 576
rect 11586 516 11590 572
rect 11590 516 11646 572
rect 11646 516 11650 572
rect 11586 512 11650 516
rect 11666 572 11730 576
rect 11666 516 11670 572
rect 11670 516 11726 572
rect 11726 516 11730 572
rect 11666 512 11730 516
rect 11746 572 11810 576
rect 11746 516 11750 572
rect 11750 516 11806 572
rect 11806 516 11810 572
rect 11746 512 11810 516
rect 15208 572 15272 576
rect 15208 516 15212 572
rect 15212 516 15268 572
rect 15268 516 15272 572
rect 15208 512 15272 516
rect 15288 572 15352 576
rect 15288 516 15292 572
rect 15292 516 15348 572
rect 15348 516 15352 572
rect 15288 512 15352 516
rect 15368 572 15432 576
rect 15368 516 15372 572
rect 15372 516 15428 572
rect 15428 516 15432 572
rect 15368 512 15432 516
rect 15448 572 15512 576
rect 15448 516 15452 572
rect 15452 516 15508 572
rect 15508 516 15512 572
rect 15448 512 15512 516
<< metal4 >>
rect 2243 15264 2563 15280
rect 2243 15200 2251 15264
rect 2315 15200 2331 15264
rect 2395 15200 2411 15264
rect 2475 15200 2491 15264
rect 2555 15200 2563 15264
rect 2243 14176 2563 15200
rect 2243 14112 2251 14176
rect 2315 14112 2331 14176
rect 2395 14112 2411 14176
rect 2475 14112 2491 14176
rect 2555 14112 2563 14176
rect 2243 13088 2563 14112
rect 2243 13024 2251 13088
rect 2315 13024 2331 13088
rect 2395 13024 2411 13088
rect 2475 13024 2491 13088
rect 2555 13024 2563 13088
rect 2243 12000 2563 13024
rect 2243 11936 2251 12000
rect 2315 11936 2331 12000
rect 2395 11936 2411 12000
rect 2475 11936 2491 12000
rect 2555 11936 2563 12000
rect 2243 10912 2563 11936
rect 2243 10848 2251 10912
rect 2315 10848 2331 10912
rect 2395 10848 2411 10912
rect 2475 10848 2491 10912
rect 2555 10848 2563 10912
rect 2243 9824 2563 10848
rect 2243 9760 2251 9824
rect 2315 9760 2331 9824
rect 2395 9760 2411 9824
rect 2475 9760 2491 9824
rect 2555 9760 2563 9824
rect 2243 8736 2563 9760
rect 2243 8672 2251 8736
rect 2315 8672 2331 8736
rect 2395 8672 2411 8736
rect 2475 8672 2491 8736
rect 2555 8672 2563 8736
rect 2243 7648 2563 8672
rect 2243 7584 2251 7648
rect 2315 7584 2331 7648
rect 2395 7584 2411 7648
rect 2475 7584 2491 7648
rect 2555 7584 2563 7648
rect 2243 6560 2563 7584
rect 2243 6496 2251 6560
rect 2315 6496 2331 6560
rect 2395 6496 2411 6560
rect 2475 6496 2491 6560
rect 2555 6496 2563 6560
rect 2243 5472 2563 6496
rect 2243 5408 2251 5472
rect 2315 5408 2331 5472
rect 2395 5408 2411 5472
rect 2475 5408 2491 5472
rect 2555 5408 2563 5472
rect 2243 4384 2563 5408
rect 2243 4320 2251 4384
rect 2315 4320 2331 4384
rect 2395 4320 2411 4384
rect 2475 4320 2491 4384
rect 2555 4320 2563 4384
rect 2243 3296 2563 4320
rect 2243 3232 2251 3296
rect 2315 3232 2331 3296
rect 2395 3232 2411 3296
rect 2475 3232 2491 3296
rect 2555 3232 2563 3296
rect 2243 2208 2563 3232
rect 2243 2144 2251 2208
rect 2315 2144 2331 2208
rect 2395 2144 2411 2208
rect 2475 2144 2491 2208
rect 2555 2144 2563 2208
rect 2243 1120 2563 2144
rect 2243 1056 2251 1120
rect 2315 1056 2331 1120
rect 2395 1056 2411 1120
rect 2475 1056 2491 1120
rect 2555 1056 2563 1120
rect 2243 496 2563 1056
rect 4094 14720 4414 15280
rect 4094 14656 4102 14720
rect 4166 14656 4182 14720
rect 4246 14656 4262 14720
rect 4326 14656 4342 14720
rect 4406 14656 4414 14720
rect 4094 13632 4414 14656
rect 4094 13568 4102 13632
rect 4166 13568 4182 13632
rect 4246 13568 4262 13632
rect 4326 13568 4342 13632
rect 4406 13568 4414 13632
rect 4094 12544 4414 13568
rect 4094 12480 4102 12544
rect 4166 12480 4182 12544
rect 4246 12480 4262 12544
rect 4326 12480 4342 12544
rect 4406 12480 4414 12544
rect 4094 11456 4414 12480
rect 4094 11392 4102 11456
rect 4166 11392 4182 11456
rect 4246 11392 4262 11456
rect 4326 11392 4342 11456
rect 4406 11392 4414 11456
rect 4094 10368 4414 11392
rect 4094 10304 4102 10368
rect 4166 10304 4182 10368
rect 4246 10304 4262 10368
rect 4326 10304 4342 10368
rect 4406 10304 4414 10368
rect 4094 9280 4414 10304
rect 4094 9216 4102 9280
rect 4166 9216 4182 9280
rect 4246 9216 4262 9280
rect 4326 9216 4342 9280
rect 4406 9216 4414 9280
rect 4094 8192 4414 9216
rect 4094 8128 4102 8192
rect 4166 8128 4182 8192
rect 4246 8128 4262 8192
rect 4326 8128 4342 8192
rect 4406 8128 4414 8192
rect 4094 7104 4414 8128
rect 4094 7040 4102 7104
rect 4166 7040 4182 7104
rect 4246 7040 4262 7104
rect 4326 7040 4342 7104
rect 4406 7040 4414 7104
rect 4094 6016 4414 7040
rect 4094 5952 4102 6016
rect 4166 5952 4182 6016
rect 4246 5952 4262 6016
rect 4326 5952 4342 6016
rect 4406 5952 4414 6016
rect 4094 4928 4414 5952
rect 4094 4864 4102 4928
rect 4166 4864 4182 4928
rect 4246 4864 4262 4928
rect 4326 4864 4342 4928
rect 4406 4864 4414 4928
rect 4094 3840 4414 4864
rect 4094 3776 4102 3840
rect 4166 3776 4182 3840
rect 4246 3776 4262 3840
rect 4326 3776 4342 3840
rect 4406 3776 4414 3840
rect 4094 2752 4414 3776
rect 4094 2688 4102 2752
rect 4166 2688 4182 2752
rect 4246 2688 4262 2752
rect 4326 2688 4342 2752
rect 4406 2688 4414 2752
rect 4094 1664 4414 2688
rect 4094 1600 4102 1664
rect 4166 1600 4182 1664
rect 4246 1600 4262 1664
rect 4326 1600 4342 1664
rect 4406 1600 4414 1664
rect 4094 576 4414 1600
rect 4094 512 4102 576
rect 4166 512 4182 576
rect 4246 512 4262 576
rect 4326 512 4342 576
rect 4406 512 4414 576
rect 4094 496 4414 512
rect 5945 15264 6265 15280
rect 5945 15200 5953 15264
rect 6017 15200 6033 15264
rect 6097 15200 6113 15264
rect 6177 15200 6193 15264
rect 6257 15200 6265 15264
rect 5945 14176 6265 15200
rect 5945 14112 5953 14176
rect 6017 14112 6033 14176
rect 6097 14112 6113 14176
rect 6177 14112 6193 14176
rect 6257 14112 6265 14176
rect 5945 13088 6265 14112
rect 5945 13024 5953 13088
rect 6017 13024 6033 13088
rect 6097 13024 6113 13088
rect 6177 13024 6193 13088
rect 6257 13024 6265 13088
rect 5945 12000 6265 13024
rect 5945 11936 5953 12000
rect 6017 11936 6033 12000
rect 6097 11936 6113 12000
rect 6177 11936 6193 12000
rect 6257 11936 6265 12000
rect 5945 10912 6265 11936
rect 5945 10848 5953 10912
rect 6017 10848 6033 10912
rect 6097 10848 6113 10912
rect 6177 10848 6193 10912
rect 6257 10848 6265 10912
rect 5945 9824 6265 10848
rect 5945 9760 5953 9824
rect 6017 9760 6033 9824
rect 6097 9760 6113 9824
rect 6177 9760 6193 9824
rect 6257 9760 6265 9824
rect 5945 8736 6265 9760
rect 5945 8672 5953 8736
rect 6017 8672 6033 8736
rect 6097 8672 6113 8736
rect 6177 8672 6193 8736
rect 6257 8672 6265 8736
rect 5945 7648 6265 8672
rect 5945 7584 5953 7648
rect 6017 7584 6033 7648
rect 6097 7584 6113 7648
rect 6177 7584 6193 7648
rect 6257 7584 6265 7648
rect 5945 6560 6265 7584
rect 5945 6496 5953 6560
rect 6017 6496 6033 6560
rect 6097 6496 6113 6560
rect 6177 6496 6193 6560
rect 6257 6496 6265 6560
rect 5945 5472 6265 6496
rect 5945 5408 5953 5472
rect 6017 5408 6033 5472
rect 6097 5408 6113 5472
rect 6177 5408 6193 5472
rect 6257 5408 6265 5472
rect 5945 4384 6265 5408
rect 5945 4320 5953 4384
rect 6017 4320 6033 4384
rect 6097 4320 6113 4384
rect 6177 4320 6193 4384
rect 6257 4320 6265 4384
rect 5945 3296 6265 4320
rect 5945 3232 5953 3296
rect 6017 3232 6033 3296
rect 6097 3232 6113 3296
rect 6177 3232 6193 3296
rect 6257 3232 6265 3296
rect 5945 2208 6265 3232
rect 5945 2144 5953 2208
rect 6017 2144 6033 2208
rect 6097 2144 6113 2208
rect 6177 2144 6193 2208
rect 6257 2144 6265 2208
rect 5945 1120 6265 2144
rect 5945 1056 5953 1120
rect 6017 1056 6033 1120
rect 6097 1056 6113 1120
rect 6177 1056 6193 1120
rect 6257 1056 6265 1120
rect 5945 496 6265 1056
rect 7796 14720 8116 15280
rect 7796 14656 7804 14720
rect 7868 14656 7884 14720
rect 7948 14656 7964 14720
rect 8028 14656 8044 14720
rect 8108 14656 8116 14720
rect 7796 13632 8116 14656
rect 7796 13568 7804 13632
rect 7868 13568 7884 13632
rect 7948 13568 7964 13632
rect 8028 13568 8044 13632
rect 8108 13568 8116 13632
rect 7796 12544 8116 13568
rect 7796 12480 7804 12544
rect 7868 12480 7884 12544
rect 7948 12480 7964 12544
rect 8028 12480 8044 12544
rect 8108 12480 8116 12544
rect 7796 11456 8116 12480
rect 7796 11392 7804 11456
rect 7868 11392 7884 11456
rect 7948 11392 7964 11456
rect 8028 11392 8044 11456
rect 8108 11392 8116 11456
rect 7796 10368 8116 11392
rect 7796 10304 7804 10368
rect 7868 10304 7884 10368
rect 7948 10304 7964 10368
rect 8028 10304 8044 10368
rect 8108 10304 8116 10368
rect 7796 9280 8116 10304
rect 7796 9216 7804 9280
rect 7868 9216 7884 9280
rect 7948 9216 7964 9280
rect 8028 9216 8044 9280
rect 8108 9216 8116 9280
rect 7796 8192 8116 9216
rect 7796 8128 7804 8192
rect 7868 8128 7884 8192
rect 7948 8128 7964 8192
rect 8028 8128 8044 8192
rect 8108 8128 8116 8192
rect 7796 7104 8116 8128
rect 7796 7040 7804 7104
rect 7868 7040 7884 7104
rect 7948 7040 7964 7104
rect 8028 7040 8044 7104
rect 8108 7040 8116 7104
rect 7796 6016 8116 7040
rect 7796 5952 7804 6016
rect 7868 5952 7884 6016
rect 7948 5952 7964 6016
rect 8028 5952 8044 6016
rect 8108 5952 8116 6016
rect 7796 4928 8116 5952
rect 7796 4864 7804 4928
rect 7868 4864 7884 4928
rect 7948 4864 7964 4928
rect 8028 4864 8044 4928
rect 8108 4864 8116 4928
rect 7796 3840 8116 4864
rect 7796 3776 7804 3840
rect 7868 3776 7884 3840
rect 7948 3776 7964 3840
rect 8028 3776 8044 3840
rect 8108 3776 8116 3840
rect 7796 2752 8116 3776
rect 7796 2688 7804 2752
rect 7868 2688 7884 2752
rect 7948 2688 7964 2752
rect 8028 2688 8044 2752
rect 8108 2688 8116 2752
rect 7796 1664 8116 2688
rect 7796 1600 7804 1664
rect 7868 1600 7884 1664
rect 7948 1600 7964 1664
rect 8028 1600 8044 1664
rect 8108 1600 8116 1664
rect 7796 576 8116 1600
rect 7796 512 7804 576
rect 7868 512 7884 576
rect 7948 512 7964 576
rect 8028 512 8044 576
rect 8108 512 8116 576
rect 7796 496 8116 512
rect 9647 15264 9967 15280
rect 9647 15200 9655 15264
rect 9719 15200 9735 15264
rect 9799 15200 9815 15264
rect 9879 15200 9895 15264
rect 9959 15200 9967 15264
rect 9647 14176 9967 15200
rect 9647 14112 9655 14176
rect 9719 14112 9735 14176
rect 9799 14112 9815 14176
rect 9879 14112 9895 14176
rect 9959 14112 9967 14176
rect 9647 13088 9967 14112
rect 9647 13024 9655 13088
rect 9719 13024 9735 13088
rect 9799 13024 9815 13088
rect 9879 13024 9895 13088
rect 9959 13024 9967 13088
rect 9647 12000 9967 13024
rect 9647 11936 9655 12000
rect 9719 11936 9735 12000
rect 9799 11936 9815 12000
rect 9879 11936 9895 12000
rect 9959 11936 9967 12000
rect 9647 10912 9967 11936
rect 9647 10848 9655 10912
rect 9719 10848 9735 10912
rect 9799 10848 9815 10912
rect 9879 10848 9895 10912
rect 9959 10848 9967 10912
rect 9647 9824 9967 10848
rect 9647 9760 9655 9824
rect 9719 9760 9735 9824
rect 9799 9760 9815 9824
rect 9879 9760 9895 9824
rect 9959 9760 9967 9824
rect 9647 8736 9967 9760
rect 9647 8672 9655 8736
rect 9719 8672 9735 8736
rect 9799 8672 9815 8736
rect 9879 8672 9895 8736
rect 9959 8672 9967 8736
rect 9647 7648 9967 8672
rect 9647 7584 9655 7648
rect 9719 7584 9735 7648
rect 9799 7584 9815 7648
rect 9879 7584 9895 7648
rect 9959 7584 9967 7648
rect 9647 6560 9967 7584
rect 9647 6496 9655 6560
rect 9719 6496 9735 6560
rect 9799 6496 9815 6560
rect 9879 6496 9895 6560
rect 9959 6496 9967 6560
rect 9647 5472 9967 6496
rect 9647 5408 9655 5472
rect 9719 5408 9735 5472
rect 9799 5408 9815 5472
rect 9879 5408 9895 5472
rect 9959 5408 9967 5472
rect 9647 4384 9967 5408
rect 9647 4320 9655 4384
rect 9719 4320 9735 4384
rect 9799 4320 9815 4384
rect 9879 4320 9895 4384
rect 9959 4320 9967 4384
rect 9647 3296 9967 4320
rect 9647 3232 9655 3296
rect 9719 3232 9735 3296
rect 9799 3232 9815 3296
rect 9879 3232 9895 3296
rect 9959 3232 9967 3296
rect 9647 2208 9967 3232
rect 9647 2144 9655 2208
rect 9719 2144 9735 2208
rect 9799 2144 9815 2208
rect 9879 2144 9895 2208
rect 9959 2144 9967 2208
rect 9647 1120 9967 2144
rect 9647 1056 9655 1120
rect 9719 1056 9735 1120
rect 9799 1056 9815 1120
rect 9879 1056 9895 1120
rect 9959 1056 9967 1120
rect 9647 496 9967 1056
rect 11498 14720 11818 15280
rect 11498 14656 11506 14720
rect 11570 14656 11586 14720
rect 11650 14656 11666 14720
rect 11730 14656 11746 14720
rect 11810 14656 11818 14720
rect 11498 13632 11818 14656
rect 11498 13568 11506 13632
rect 11570 13568 11586 13632
rect 11650 13568 11666 13632
rect 11730 13568 11746 13632
rect 11810 13568 11818 13632
rect 11498 12544 11818 13568
rect 11498 12480 11506 12544
rect 11570 12480 11586 12544
rect 11650 12480 11666 12544
rect 11730 12480 11746 12544
rect 11810 12480 11818 12544
rect 11498 11456 11818 12480
rect 11498 11392 11506 11456
rect 11570 11392 11586 11456
rect 11650 11392 11666 11456
rect 11730 11392 11746 11456
rect 11810 11392 11818 11456
rect 11498 10368 11818 11392
rect 11498 10304 11506 10368
rect 11570 10304 11586 10368
rect 11650 10304 11666 10368
rect 11730 10304 11746 10368
rect 11810 10304 11818 10368
rect 11498 9280 11818 10304
rect 11498 9216 11506 9280
rect 11570 9216 11586 9280
rect 11650 9216 11666 9280
rect 11730 9216 11746 9280
rect 11810 9216 11818 9280
rect 11498 8192 11818 9216
rect 11498 8128 11506 8192
rect 11570 8128 11586 8192
rect 11650 8128 11666 8192
rect 11730 8128 11746 8192
rect 11810 8128 11818 8192
rect 11498 7104 11818 8128
rect 11498 7040 11506 7104
rect 11570 7040 11586 7104
rect 11650 7040 11666 7104
rect 11730 7040 11746 7104
rect 11810 7040 11818 7104
rect 11498 6016 11818 7040
rect 11498 5952 11506 6016
rect 11570 5952 11586 6016
rect 11650 5952 11666 6016
rect 11730 5952 11746 6016
rect 11810 5952 11818 6016
rect 11498 4928 11818 5952
rect 11498 4864 11506 4928
rect 11570 4864 11586 4928
rect 11650 4864 11666 4928
rect 11730 4864 11746 4928
rect 11810 4864 11818 4928
rect 11498 3840 11818 4864
rect 11498 3776 11506 3840
rect 11570 3776 11586 3840
rect 11650 3776 11666 3840
rect 11730 3776 11746 3840
rect 11810 3776 11818 3840
rect 11498 2752 11818 3776
rect 11498 2688 11506 2752
rect 11570 2688 11586 2752
rect 11650 2688 11666 2752
rect 11730 2688 11746 2752
rect 11810 2688 11818 2752
rect 11498 1664 11818 2688
rect 11498 1600 11506 1664
rect 11570 1600 11586 1664
rect 11650 1600 11666 1664
rect 11730 1600 11746 1664
rect 11810 1600 11818 1664
rect 11498 576 11818 1600
rect 11498 512 11506 576
rect 11570 512 11586 576
rect 11650 512 11666 576
rect 11730 512 11746 576
rect 11810 512 11818 576
rect 11498 496 11818 512
rect 13349 15264 13669 15280
rect 13349 15200 13357 15264
rect 13421 15200 13437 15264
rect 13501 15200 13517 15264
rect 13581 15200 13597 15264
rect 13661 15200 13669 15264
rect 13349 14176 13669 15200
rect 13349 14112 13357 14176
rect 13421 14112 13437 14176
rect 13501 14112 13517 14176
rect 13581 14112 13597 14176
rect 13661 14112 13669 14176
rect 13349 13088 13669 14112
rect 13349 13024 13357 13088
rect 13421 13024 13437 13088
rect 13501 13024 13517 13088
rect 13581 13024 13597 13088
rect 13661 13024 13669 13088
rect 13349 12000 13669 13024
rect 13349 11936 13357 12000
rect 13421 11936 13437 12000
rect 13501 11936 13517 12000
rect 13581 11936 13597 12000
rect 13661 11936 13669 12000
rect 13349 10912 13669 11936
rect 13349 10848 13357 10912
rect 13421 10848 13437 10912
rect 13501 10848 13517 10912
rect 13581 10848 13597 10912
rect 13661 10848 13669 10912
rect 13349 9824 13669 10848
rect 13349 9760 13357 9824
rect 13421 9760 13437 9824
rect 13501 9760 13517 9824
rect 13581 9760 13597 9824
rect 13661 9760 13669 9824
rect 13349 8736 13669 9760
rect 13349 8672 13357 8736
rect 13421 8672 13437 8736
rect 13501 8672 13517 8736
rect 13581 8672 13597 8736
rect 13661 8672 13669 8736
rect 13349 7648 13669 8672
rect 13349 7584 13357 7648
rect 13421 7584 13437 7648
rect 13501 7584 13517 7648
rect 13581 7584 13597 7648
rect 13661 7584 13669 7648
rect 13349 6560 13669 7584
rect 13349 6496 13357 6560
rect 13421 6496 13437 6560
rect 13501 6496 13517 6560
rect 13581 6496 13597 6560
rect 13661 6496 13669 6560
rect 13349 5472 13669 6496
rect 13349 5408 13357 5472
rect 13421 5408 13437 5472
rect 13501 5408 13517 5472
rect 13581 5408 13597 5472
rect 13661 5408 13669 5472
rect 13349 4384 13669 5408
rect 13349 4320 13357 4384
rect 13421 4320 13437 4384
rect 13501 4320 13517 4384
rect 13581 4320 13597 4384
rect 13661 4320 13669 4384
rect 13349 3296 13669 4320
rect 13349 3232 13357 3296
rect 13421 3232 13437 3296
rect 13501 3232 13517 3296
rect 13581 3232 13597 3296
rect 13661 3232 13669 3296
rect 13349 2208 13669 3232
rect 13349 2144 13357 2208
rect 13421 2144 13437 2208
rect 13501 2144 13517 2208
rect 13581 2144 13597 2208
rect 13661 2144 13669 2208
rect 13349 1120 13669 2144
rect 13349 1056 13357 1120
rect 13421 1056 13437 1120
rect 13501 1056 13517 1120
rect 13581 1056 13597 1120
rect 13661 1056 13669 1120
rect 13349 496 13669 1056
rect 15200 14720 15520 15280
rect 15200 14656 15208 14720
rect 15272 14656 15288 14720
rect 15352 14656 15368 14720
rect 15432 14656 15448 14720
rect 15512 14656 15520 14720
rect 15200 13632 15520 14656
rect 15200 13568 15208 13632
rect 15272 13568 15288 13632
rect 15352 13568 15368 13632
rect 15432 13568 15448 13632
rect 15512 13568 15520 13632
rect 15200 12544 15520 13568
rect 15200 12480 15208 12544
rect 15272 12480 15288 12544
rect 15352 12480 15368 12544
rect 15432 12480 15448 12544
rect 15512 12480 15520 12544
rect 15200 11456 15520 12480
rect 15200 11392 15208 11456
rect 15272 11392 15288 11456
rect 15352 11392 15368 11456
rect 15432 11392 15448 11456
rect 15512 11392 15520 11456
rect 15200 10368 15520 11392
rect 15200 10304 15208 10368
rect 15272 10304 15288 10368
rect 15352 10304 15368 10368
rect 15432 10304 15448 10368
rect 15512 10304 15520 10368
rect 15200 9280 15520 10304
rect 15200 9216 15208 9280
rect 15272 9216 15288 9280
rect 15352 9216 15368 9280
rect 15432 9216 15448 9280
rect 15512 9216 15520 9280
rect 15200 8192 15520 9216
rect 15200 8128 15208 8192
rect 15272 8128 15288 8192
rect 15352 8128 15368 8192
rect 15432 8128 15448 8192
rect 15512 8128 15520 8192
rect 15200 7104 15520 8128
rect 15200 7040 15208 7104
rect 15272 7040 15288 7104
rect 15352 7040 15368 7104
rect 15432 7040 15448 7104
rect 15512 7040 15520 7104
rect 15200 6016 15520 7040
rect 15200 5952 15208 6016
rect 15272 5952 15288 6016
rect 15352 5952 15368 6016
rect 15432 5952 15448 6016
rect 15512 5952 15520 6016
rect 15200 4928 15520 5952
rect 15200 4864 15208 4928
rect 15272 4864 15288 4928
rect 15352 4864 15368 4928
rect 15432 4864 15448 4928
rect 15512 4864 15520 4928
rect 15200 3840 15520 4864
rect 15200 3776 15208 3840
rect 15272 3776 15288 3840
rect 15352 3776 15368 3840
rect 15432 3776 15448 3840
rect 15512 3776 15520 3840
rect 15200 2752 15520 3776
rect 15200 2688 15208 2752
rect 15272 2688 15288 2752
rect 15352 2688 15368 2752
rect 15432 2688 15448 2752
rect 15512 2688 15520 2752
rect 15200 1664 15520 2688
rect 15200 1600 15208 1664
rect 15272 1600 15288 1664
rect 15352 1600 15368 1664
rect 15432 1600 15448 1664
rect 15512 1600 15520 1664
rect 15200 576 15520 1600
rect 15200 512 15208 576
rect 15272 512 15288 576
rect 15352 512 15368 576
rect 15432 512 15448 576
rect 15512 512 15520 576
rect 15200 496 15520 512
use sky130_fd_sc_hd__nand2_1  _048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 6992 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_2  _049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8648 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7176 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7728 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__a41o_1  _055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5980 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _056_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5336 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _057_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7912 0 1 11424
box -38 -48 498 592
use sky130_fd_sc_hd__o22ai_1  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5244 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _059_
timestamp 1704896540
transform -1 0 8832 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _060_
timestamp 1704896540
transform -1 0 5704 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7728 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__and3b_1  _062_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7176 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__nand2b_2  _064_
timestamp 1704896540
transform 1 0 8924 0 1 11424
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _065_
timestamp 1704896540
transform -1 0 10580 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10120 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8556 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _068_
timestamp 1704896540
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _069_
timestamp 1704896540
transform 1 0 9660 0 -1 13600
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _070_
timestamp 1704896540
transform 1 0 12788 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _071_
timestamp 1704896540
transform 1 0 10672 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _072_
timestamp 1704896540
transform -1 0 10764 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _073_
timestamp 1704896540
transform 1 0 9936 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 13600
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _075_
timestamp 1704896540
transform -1 0 8924 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _076_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9200 0 -1 12512
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _077_
timestamp 1704896540
transform 1 0 12696 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _078_
timestamp 1704896540
transform 1 0 12144 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _079_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 10764 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9384 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _081_
timestamp 1704896540
transform -1 0 10672 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _082_
timestamp 1704896540
transform 1 0 6256 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8832 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _084_
timestamp 1704896540
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _085_
timestamp 1704896540
transform 1 0 14444 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _086_
timestamp 1704896540
transform 1 0 8464 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _087_
timestamp 1704896540
transform 1 0 6440 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _088_
timestamp 1704896540
transform -1 0 6348 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _089_
timestamp 1704896540
transform -1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _090_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4600 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1704896540
transform -1 0 10396 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1704896540
transform -1 0 8280 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 1704896540
transform 1 0 6716 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1704896540
transform 1 0 11408 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1704896540
transform 1 0 12512 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1704896540
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1704896540
transform -1 0 10856 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1704896540
transform 1 0 7728 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1704896540
transform -1 0 6072 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1704896540
transform -1 0 6072 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1704896540
transform 1 0 4600 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1704896540
transform -1 0 3956 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _103_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9108 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_2  _104_
timestamp 1704896540
transform -1 0 9200 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _105_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5796 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _106_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10948 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _107_
timestamp 1704896540
transform 1 0 10948 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _108_
timestamp 1704896540
transform 1 0 10948 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _109_
timestamp 1704896540
transform 1 0 8740 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _110_
timestamp 1704896540
transform 1 0 6716 0 -1 14688
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _111_
timestamp 1704896540
transform 1 0 4600 0 1 13600
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _112_
timestamp 1704896540
transform 1 0 3864 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _113_
timestamp 1704896540
transform 1 0 3864 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__conb_1  _114__3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _114_
timestamp 1704896540
transform 1 0 2024 0 -1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6440 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704896540
transform -1 0 6348 0 1 12512
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704896540
transform 1 0 9568 0 1 11424
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 828 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 1932 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1704896540
transform 1 0 3220 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1704896540
transform 1 0 4324 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704896540
transform 1 0 5796 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1704896540
transform 1 0 6900 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1704896540
transform 1 0 8004 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_89
timestamp 1704896540
transform 1 0 8740 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_101 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9844 0 1 544
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1704896540
transform 1 0 10580 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1704896540
transform 1 0 10948 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1704896540
transform 1 0 12052 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1704896540
transform 1 0 13156 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1704896540
transform 1 0 13524 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_153 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 14628 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_157
timestamp 1704896540
transform 1 0 14996 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 828 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 1932 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3036 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1704896540
transform 1 0 4140 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1704896540
transform 1 0 5244 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704896540
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1704896540
transform 1 0 5796 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1704896540
transform 1 0 6900 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1704896540
transform 1 0 8004 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1704896540
transform 1 0 9108 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10212 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1704896540
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1704896540
transform 1 0 10948 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1704896540
transform 1 0 12052 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1704896540
transform 1 0 13156 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_149
timestamp 1704896540
transform 1 0 14260 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_157
timestamp 1704896540
transform 1 0 14996 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 828 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 1932 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3220 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1704896540
transform 1 0 4324 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1704896540
transform 1 0 5428 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1704896540
transform 1 0 6532 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1704896540
transform 1 0 7636 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1704896540
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1704896540
transform 1 0 8372 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1704896540
transform 1 0 9476 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1704896540
transform 1 0 10580 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1704896540
transform 1 0 11684 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1704896540
transform 1 0 12788 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1704896540
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1704896540
transform 1 0 13524 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 1704896540
transform 1 0 14628 0 1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1704896540
transform 1 0 14996 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 828 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 1932 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3036 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4140 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1704896540
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1704896540
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704896540
transform 1 0 5796 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1704896540
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1704896540
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1704896540
transform 1 0 9108 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1704896540
transform 1 0 10212 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1704896540
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1704896540
transform 1 0 10948 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1704896540
transform 1 0 12052 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1704896540
transform 1 0 13156 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_149
timestamp 1704896540
transform 1 0 14260 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_157
timestamp 1704896540
transform 1 0 14996 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 828 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 1932 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3220 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4324 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1704896540
transform 1 0 5428 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1704896540
transform 1 0 6532 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1704896540
transform 1 0 7636 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8372 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1704896540
transform 1 0 9476 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1704896540
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1704896540
transform 1 0 11684 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1704896540
transform 1 0 12788 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1704896540
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1704896540
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_153
timestamp 1704896540
transform 1 0 14628 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_157
timestamp 1704896540
transform 1 0 14996 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 828 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1704896540
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1704896540
transform 1 0 3036 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1704896540
transform 1 0 4140 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1704896540
transform 1 0 5244 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1704896540
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1704896540
transform 1 0 5796 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1704896540
transform 1 0 6900 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1704896540
transform 1 0 8004 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1704896540
transform 1 0 9108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1704896540
transform 1 0 10212 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1704896540
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1704896540
transform 1 0 10948 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1704896540
transform 1 0 12052 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1704896540
transform 1 0 13156 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_149
timestamp 1704896540
transform 1 0 14260 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_157
timestamp 1704896540
transform 1 0 14996 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 828 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1704896540
transform 1 0 1932 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1704896540
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1704896540
transform 1 0 3220 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1704896540
transform 1 0 4324 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1704896540
transform 1 0 5428 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1704896540
transform 1 0 6532 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1704896540
transform 1 0 7636 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1704896540
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1704896540
transform 1 0 8372 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1704896540
transform 1 0 9476 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1704896540
transform 1 0 10580 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1704896540
transform 1 0 11684 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1704896540
transform 1 0 12788 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1704896540
transform 1 0 13340 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1704896540
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 1704896540
transform 1 0 14628 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1704896540
transform 1 0 14996 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 828 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 1932 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3036 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4140 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1704896540
transform 1 0 5244 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1704896540
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1704896540
transform 1 0 5796 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1704896540
transform 1 0 6900 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1704896540
transform 1 0 8004 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1704896540
transform 1 0 9108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1704896540
transform 1 0 10212 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1704896540
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1704896540
transform 1 0 10948 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1704896540
transform 1 0 12052 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1704896540
transform 1 0 13156 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_149
timestamp 1704896540
transform 1 0 14260 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_157
timestamp 1704896540
transform 1 0 14996 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1704896540
transform 1 0 828 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1704896540
transform 1 0 1932 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1704896540
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3220 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1704896540
transform 1 0 4324 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1704896540
transform 1 0 5428 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1704896540
transform 1 0 6532 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1704896540
transform 1 0 7636 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1704896540
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8372 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1704896540
transform 1 0 9476 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1704896540
transform 1 0 10580 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1704896540
transform 1 0 11684 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1704896540
transform 1 0 12788 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1704896540
transform 1 0 13340 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1704896540
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_153
timestamp 1704896540
transform 1 0 14628 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_157
timestamp 1704896540
transform 1 0 14996 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 828 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1704896540
transform 1 0 1932 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3036 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1704896540
transform 1 0 4140 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1704896540
transform 1 0 5244 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1704896540
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1704896540
transform 1 0 5796 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1704896540
transform 1 0 6900 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1704896540
transform 1 0 8004 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1704896540
transform 1 0 9108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1704896540
transform 1 0 10212 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1704896540
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1704896540
transform 1 0 10948 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1704896540
transform 1 0 12052 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1704896540
transform 1 0 13156 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_149
timestamp 1704896540
transform 1 0 14260 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_157
timestamp 1704896540
transform 1 0 14996 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 828 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 1932 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3220 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4324 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1704896540
transform 1 0 5428 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1704896540
transform 1 0 6532 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1704896540
transform 1 0 7636 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1704896540
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8372 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1704896540
transform 1 0 9476 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1704896540
transform 1 0 10580 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1704896540
transform 1 0 11684 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1704896540
transform 1 0 12788 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1704896540
transform 1 0 13340 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1704896540
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_153
timestamp 1704896540
transform 1 0 14628 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_157
timestamp 1704896540
transform 1 0 14996 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 828 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1704896540
transform 1 0 1932 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3036 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1704896540
transform 1 0 4140 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1704896540
transform 1 0 5244 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1704896540
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1704896540
transform 1 0 5796 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1704896540
transform 1 0 6900 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1704896540
transform 1 0 8004 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1704896540
transform 1 0 9108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1704896540
transform 1 0 10212 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1704896540
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1704896540
transform 1 0 10948 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1704896540
transform 1 0 12052 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13156 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_149
timestamp 1704896540
transform 1 0 14260 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_157
timestamp 1704896540
transform 1 0 14996 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1704896540
transform 1 0 828 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1704896540
transform 1 0 1932 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3220 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1704896540
transform 1 0 4324 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1704896540
transform 1 0 5428 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1704896540
transform 1 0 6532 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1704896540
transform 1 0 7636 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1704896540
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1704896540
transform 1 0 8372 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1704896540
transform 1 0 9476 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1704896540
transform 1 0 10580 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1704896540
transform 1 0 11684 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1704896540
transform 1 0 12788 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13340 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1704896540
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_153
timestamp 1704896540
transform 1 0 14628 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_157
timestamp 1704896540
transform 1 0 14996 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704896540
transform 1 0 828 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704896540
transform 1 0 1932 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1704896540
transform 1 0 3036 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1704896540
transform 1 0 4140 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1704896540
transform 1 0 5244 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1704896540
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1704896540
transform 1 0 5796 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1704896540
transform 1 0 6900 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1704896540
transform 1 0 8004 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1704896540
transform 1 0 10212 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1704896540
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1704896540
transform 1 0 10948 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1704896540
transform 1 0 12052 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1704896540
transform 1 0 13156 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_149
timestamp 1704896540
transform 1 0 14260 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_157
timestamp 1704896540
transform 1 0 14996 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1704896540
transform 1 0 828 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1704896540
transform 1 0 1932 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3220 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4324 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5428 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1704896540
transform 1 0 6532 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1704896540
transform 1 0 7636 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1704896540
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8372 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1704896540
transform 1 0 9476 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1704896540
transform 1 0 10580 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1704896540
transform 1 0 11684 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1704896540
transform 1 0 12788 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1704896540
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1704896540
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1704896540
transform 1 0 14628 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1704896540
transform 1 0 14996 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1704896540
transform 1 0 828 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1704896540
transform 1 0 1932 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1704896540
transform 1 0 3036 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1704896540
transform 1 0 4140 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1704896540
transform 1 0 5244 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1704896540
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1704896540
transform 1 0 5796 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1704896540
transform 1 0 6900 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1704896540
transform 1 0 8004 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1704896540
transform 1 0 9108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1704896540
transform 1 0 10212 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1704896540
transform 1 0 10948 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1704896540
transform 1 0 12052 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1704896540
transform 1 0 13156 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_149
timestamp 1704896540
transform 1 0 14260 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_157
timestamp 1704896540
transform 1 0 14996 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1704896540
transform 1 0 828 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1704896540
transform 1 0 1932 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1704896540
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1704896540
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_53
timestamp 1704896540
transform 1 0 5428 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_61
timestamp 1704896540
transform 1 0 6164 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_68
timestamp 1704896540
transform 1 0 6808 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_80
timestamp 1704896540
transform 1 0 7912 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8372 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1704896540
transform 1 0 9476 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1704896540
transform 1 0 10580 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1704896540
transform 1 0 11684 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1704896540
transform 1 0 12788 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1704896540
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1704896540
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_153
timestamp 1704896540
transform 1 0 14628 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_157
timestamp 1704896540
transform 1 0 14996 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1704896540
transform 1 0 828 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1704896540
transform 1 0 1932 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1704896540
transform 1 0 3036 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1704896540
transform 1 0 4140 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5244 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1704896540
transform 1 0 5796 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_61
timestamp 1704896540
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_70
timestamp 1704896540
transform 1 0 6992 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_94
timestamp 1704896540
transform 1 0 9200 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_102 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9936 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 1704896540
transform 1 0 10396 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1704896540
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1704896540
transform 1 0 10948 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1704896540
transform 1 0 12052 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1704896540
transform 1 0 13156 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_149
timestamp 1704896540
transform 1 0 14260 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_157
timestamp 1704896540
transform 1 0 14996 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1704896540
transform 1 0 828 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1704896540
transform 1 0 1932 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1704896540
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3220 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1704896540
transform 1 0 4324 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_53
timestamp 1704896540
transform 1 0 5428 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_78
timestamp 1704896540
transform 1 0 7728 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_114
timestamp 1704896540
transform 1 0 11040 0 1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1704896540
transform 1 0 11684 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1704896540
transform 1 0 12788 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1704896540
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_153
timestamp 1704896540
transform 1 0 14628 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_157
timestamp 1704896540
transform 1 0 14996 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1704896540
transform 1 0 828 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1704896540
transform 1 0 1932 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_27
timestamp 1704896540
transform 1 0 3036 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_35
timestamp 1704896540
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_60
timestamp 1704896540
transform 1 0 6072 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_66
timestamp 1704896540
transform 1 0 6624 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_70
timestamp 1704896540
transform 1 0 6992 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_90
timestamp 1704896540
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_110
timestamp 1704896540
transform 1 0 10672 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_133
timestamp 1704896540
transform 1 0 12788 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_145
timestamp 1704896540
transform 1 0 13892 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_157
timestamp 1704896540
transform 1 0 14996 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1704896540
transform 1 0 828 0 1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1704896540
transform 1 0 1932 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1704896540
transform 1 0 3036 0 1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3220 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_41
timestamp 1704896540
transform 1 0 4324 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_47
timestamp 1704896540
transform 1 0 4876 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_51
timestamp 1704896540
transform 1 0 5244 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_80
timestamp 1704896540
transform 1 0 7912 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8372 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1704896540
transform 1 0 12788 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1704896540
transform 1 0 13340 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1704896540
transform 1 0 13524 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_149
timestamp 1704896540
transform 1 0 14260 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_154
timestamp 1704896540
transform 1 0 14720 0 1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1704896540
transform 1 0 828 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_15
timestamp 1704896540
transform 1 0 1932 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_65
timestamp 1704896540
transform 1 0 6532 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_70
timestamp 1704896540
transform 1 0 6992 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_87
timestamp 1704896540
transform 1 0 8556 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_91
timestamp 1704896540
transform 1 0 8924 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_101
timestamp 1704896540
transform 1 0 9844 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1704896540
transform 1 0 10764 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_133
timestamp 1704896540
transform 1 0 12788 0 -1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_145
timestamp 1704896540
transform 1 0 13892 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_157
timestamp 1704896540
transform 1 0 14996 0 -1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1704896540
transform 1 0 828 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1704896540
transform 1 0 1932 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1704896540
transform 1 0 3036 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3220 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_63
timestamp 1704896540
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_92
timestamp 1704896540
transform 1 0 9016 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_100
timestamp 1704896540
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_105
timestamp 1704896540
transform 1 0 10212 0 1 12512
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_117
timestamp 1704896540
transform 1 0 11316 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_129
timestamp 1704896540
transform 1 0 12420 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 1704896540
transform 1 0 12972 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1704896540
transform 1 0 13340 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1704896540
transform 1 0 13524 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_153
timestamp 1704896540
transform 1 0 14628 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_157
timestamp 1704896540
transform 1 0 14996 0 1 12512
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1704896540
transform 1 0 828 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1704896540
transform 1 0 1932 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_30
timestamp 1704896540
transform 1 0 3312 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_37
timestamp 1704896540
transform 1 0 3956 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_45
timestamp 1704896540
transform 1 0 4692 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1704896540
transform 1 0 5796 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_98
timestamp 1704896540
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1704896540
transform 1 0 10764 0 -1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_120
timestamp 1704896540
transform 1 0 11592 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_132
timestamp 1704896540
transform 1 0 12696 0 -1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_144
timestamp 1704896540
transform 1 0 13800 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_156
timestamp 1704896540
transform 1 0 14904 0 -1 13600
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1704896540
transform 1 0 828 0 1 13600
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1704896540
transform 1 0 1932 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1704896540
transform 1 0 3036 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1704896540
transform 1 0 3220 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_41
timestamp 1704896540
transform 1 0 4324 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1704896540
transform 1 0 8004 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_97
timestamp 1704896540
transform 1 0 9476 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_105
timestamp 1704896540
transform 1 0 10212 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_109
timestamp 1704896540
transform 1 0 10580 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_114
timestamp 1704896540
transform 1 0 11040 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_120
timestamp 1704896540
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_124
timestamp 1704896540
transform 1 0 11960 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1704896540
transform 1 0 13064 0 1 13600
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1704896540
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_153
timestamp 1704896540
transform 1 0 14628 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_157
timestamp 1704896540
transform 1 0 14996 0 1 13600
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 828 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1704896540
transform 1 0 1932 0 -1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1704896540
transform 1 0 3036 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_39
timestamp 1704896540
transform 1 0 4140 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_43
timestamp 1704896540
transform 1 0 4508 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1704896540
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_63
timestamp 1704896540
transform 1 0 6348 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_87
timestamp 1704896540
transform 1 0 8556 0 -1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_136
timestamp 1704896540
transform 1 0 13064 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_148
timestamp 1704896540
transform 1 0 14168 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_156
timestamp 1704896540
transform 1 0 14904 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1704896540
transform 1 0 828 0 1 14688
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_8
timestamp 1704896540
transform 1 0 1288 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_20
timestamp 1704896540
transform 1 0 2392 0 1 14688
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1704896540
transform 1 0 3220 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1704896540
transform 1 0 4324 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_53
timestamp 1704896540
transform 1 0 5428 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_57
timestamp 1704896540
transform 1 0 5796 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_69
timestamp 1704896540
transform 1 0 6900 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1704896540
transform 1 0 8004 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 1704896540
transform 1 0 8372 0 1 14688
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_89
timestamp 1704896540
transform 1 0 8740 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_101
timestamp 1704896540
transform 1 0 9844 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_109
timestamp 1704896540
transform 1 0 10580 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_113
timestamp 1704896540
transform 1 0 10948 0 1 14688
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_125
timestamp 1704896540
transform 1 0 12052 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_137
timestamp 1704896540
transform 1 0 13156 0 1 14688
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 13524 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_153
timestamp 1704896540
transform 1 0 14628 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_157
timestamp 1704896540
transform 1 0 14996 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 9108 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 12144 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform 1 0 6440 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform 1 0 5980 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 9108 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 6992 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform 1 0 7544 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 7452 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 544
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1012 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_27
timestamp 1704896540
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 15364 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_28
timestamp 1704896540
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 15364 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_29
timestamp 1704896540
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 15364 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_30
timestamp 1704896540
transform 1 0 552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 15364 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_31
timestamp 1704896540
transform 1 0 552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 15364 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_32
timestamp 1704896540
transform 1 0 552 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 15364 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_33
timestamp 1704896540
transform 1 0 552 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 15364 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_34
timestamp 1704896540
transform 1 0 552 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 15364 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_35
timestamp 1704896540
transform 1 0 552 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 15364 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_36
timestamp 1704896540
transform 1 0 552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 15364 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_37
timestamp 1704896540
transform 1 0 552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 15364 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_38
timestamp 1704896540
transform 1 0 552 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 15364 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_39
timestamp 1704896540
transform 1 0 552 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 15364 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_40
timestamp 1704896540
transform 1 0 552 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 15364 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_41
timestamp 1704896540
transform 1 0 552 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 15364 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_42
timestamp 1704896540
transform 1 0 552 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 15364 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_43
timestamp 1704896540
transform 1 0 552 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 15364 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_44
timestamp 1704896540
transform 1 0 552 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 15364 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_45
timestamp 1704896540
transform 1 0 552 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 15364 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_46
timestamp 1704896540
transform 1 0 552 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 15364 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_47
timestamp 1704896540
transform 1 0 552 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 15364 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_48
timestamp 1704896540
transform 1 0 552 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 15364 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_49
timestamp 1704896540
transform 1 0 552 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 15364 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_50
timestamp 1704896540
transform 1 0 552 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 15364 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_51
timestamp 1704896540
transform 1 0 552 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 15364 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_52
timestamp 1704896540
transform 1 0 552 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 15364 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_53
timestamp 1704896540
transform 1 0 552 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 15364 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_55
timestamp 1704896540
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_56
timestamp 1704896540
transform 1 0 8280 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_57
timestamp 1704896540
transform 1 0 10856 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 1704896540
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_59
timestamp 1704896540
transform 1 0 5704 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_60
timestamp 1704896540
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_61
timestamp 1704896540
transform 1 0 3128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_62
timestamp 1704896540
transform 1 0 8280 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_63
timestamp 1704896540
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_64
timestamp 1704896540
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_65
timestamp 1704896540
transform 1 0 10856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp 1704896540
transform 1 0 3128 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp 1704896540
transform 1 0 8280 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp 1704896540
transform 1 0 13432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_69
timestamp 1704896540
transform 1 0 5704 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp 1704896540
transform 1 0 10856 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_71
timestamp 1704896540
transform 1 0 3128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_72
timestamp 1704896540
transform 1 0 8280 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_73
timestamp 1704896540
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_74
timestamp 1704896540
transform 1 0 5704 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_75
timestamp 1704896540
transform 1 0 10856 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_76
timestamp 1704896540
transform 1 0 3128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_77
timestamp 1704896540
transform 1 0 8280 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_78
timestamp 1704896540
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_79
timestamp 1704896540
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_80
timestamp 1704896540
transform 1 0 10856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_81
timestamp 1704896540
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_82
timestamp 1704896540
transform 1 0 8280 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_83
timestamp 1704896540
transform 1 0 13432 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_84
timestamp 1704896540
transform 1 0 5704 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_85
timestamp 1704896540
transform 1 0 10856 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_86
timestamp 1704896540
transform 1 0 3128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_87
timestamp 1704896540
transform 1 0 8280 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_88
timestamp 1704896540
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_89
timestamp 1704896540
transform 1 0 5704 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_90
timestamp 1704896540
transform 1 0 10856 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_91
timestamp 1704896540
transform 1 0 3128 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_92
timestamp 1704896540
transform 1 0 8280 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_93
timestamp 1704896540
transform 1 0 13432 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_94
timestamp 1704896540
transform 1 0 5704 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_95
timestamp 1704896540
transform 1 0 10856 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_96
timestamp 1704896540
transform 1 0 3128 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_97
timestamp 1704896540
transform 1 0 8280 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_98
timestamp 1704896540
transform 1 0 13432 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_99
timestamp 1704896540
transform 1 0 5704 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_100
timestamp 1704896540
transform 1 0 10856 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_101
timestamp 1704896540
transform 1 0 3128 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_102
timestamp 1704896540
transform 1 0 8280 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_103
timestamp 1704896540
transform 1 0 13432 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_104
timestamp 1704896540
transform 1 0 5704 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_105
timestamp 1704896540
transform 1 0 10856 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_106
timestamp 1704896540
transform 1 0 3128 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_107
timestamp 1704896540
transform 1 0 8280 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_108
timestamp 1704896540
transform 1 0 13432 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_109
timestamp 1704896540
transform 1 0 5704 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_110
timestamp 1704896540
transform 1 0 10856 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_111
timestamp 1704896540
transform 1 0 3128 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_112
timestamp 1704896540
transform 1 0 8280 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_113
timestamp 1704896540
transform 1 0 13432 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_114
timestamp 1704896540
transform 1 0 5704 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_115
timestamp 1704896540
transform 1 0 10856 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_116
timestamp 1704896540
transform 1 0 3128 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_117
timestamp 1704896540
transform 1 0 8280 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_118
timestamp 1704896540
transform 1 0 13432 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_119
timestamp 1704896540
transform 1 0 5704 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_120
timestamp 1704896540
transform 1 0 10856 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_121
timestamp 1704896540
transform 1 0 3128 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_122
timestamp 1704896540
transform 1 0 5704 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_123
timestamp 1704896540
transform 1 0 8280 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_124
timestamp 1704896540
transform 1 0 10856 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_125
timestamp 1704896540
transform 1 0 13432 0 1 14688
box -38 -48 130 592
<< labels >>
flabel metal4 s 4094 496 4414 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7796 496 8116 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 11498 496 11818 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 15200 496 15520 15280 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2243 496 2563 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 5945 496 6265 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 9647 496 9967 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 13349 496 13669 15280 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 2502 15600 2558 16000 0 FreeSans 224 90 0 0 clk
port 2 nsew signal input
flabel metal2 s 7930 0 7986 400 0 FreeSans 224 90 0 0 comp
port 3 nsew signal input
flabel metal2 s 15014 15600 15070 16000 0 FreeSans 224 90 0 0 data_out[0]
port 4 nsew signal output
flabel metal2 s 13450 15600 13506 16000 0 FreeSans 224 90 0 0 data_out[1]
port 5 nsew signal output
flabel metal2 s 11886 15600 11942 16000 0 FreeSans 224 90 0 0 data_out[2]
port 6 nsew signal output
flabel metal2 s 10322 15600 10378 16000 0 FreeSans 224 90 0 0 data_out[3]
port 7 nsew signal output
flabel metal2 s 8758 15600 8814 16000 0 FreeSans 224 90 0 0 data_out[4]
port 8 nsew signal output
flabel metal2 s 7194 15600 7250 16000 0 FreeSans 224 90 0 0 data_out[5]
port 9 nsew signal output
flabel metal2 s 5630 15600 5686 16000 0 FreeSans 224 90 0 0 data_out[6]
port 10 nsew signal output
flabel metal2 s 4066 15600 4122 16000 0 FreeSans 224 90 0 0 data_out[7]
port 11 nsew signal output
flabel metal2 s 938 15600 994 16000 0 FreeSans 224 90 0 0 reset
port 12 nsew signal input
rlabel via1 8036 14688 8036 14688 0 VGND
rlabel metal1 7958 15232 7958 15232 0 VPWR
rlabel metal2 10258 10370 10258 10370 0 _000_
rlabel metal2 8234 10302 8234 10302 0 _001_
rlabel metal1 6900 11050 6900 11050 0 _002_
rlabel metal2 11546 11016 11546 11016 0 _003_
rlabel metal2 12650 12070 12650 12070 0 _004_
rlabel metal2 11822 14280 11822 14280 0 _005_
rlabel metal1 10495 14518 10495 14518 0 _006_
rlabel metal1 7820 14042 7820 14042 0 _007_
rlabel metal2 5658 14008 5658 14008 0 _008_
rlabel metal1 5665 11254 5665 11254 0 _009_
rlabel metal2 4738 12104 4738 12104 0 _010_
rlabel metal1 3687 12342 3687 12342 0 _011_
rlabel metal1 9384 10574 9384 10574 0 _012_
rlabel metal2 8786 10540 8786 10540 0 _013_
rlabel metal1 6624 9622 6624 9622 0 _014_
rlabel metal1 10948 11254 10948 11254 0 _015_
rlabel metal1 10994 12342 10994 12342 0 _016_
rlabel metal1 11408 13498 11408 13498 0 _017_
rlabel metal1 8970 13498 8970 13498 0 _018_
rlabel metal1 7130 13498 7130 13498 0 _019_
rlabel metal1 6302 13872 6302 13872 0 _020_
rlabel metal1 4784 11118 4784 11118 0 _021_
rlabel metal1 5014 12206 5014 12206 0 _022_
rlabel metal1 5566 13294 5566 13294 0 _023_
rlabel metal1 5566 12954 5566 12954 0 _024_
rlabel metal1 7912 12954 7912 12954 0 _025_
rlabel metal1 6670 13226 6670 13226 0 _026_
rlabel metal1 8188 13158 8188 13158 0 _027_
rlabel metal1 5244 12818 5244 12818 0 _028_
rlabel metal1 5934 11662 5934 11662 0 _029_
rlabel metal1 5336 13158 5336 13158 0 _030_
rlabel metal1 5014 13192 5014 13192 0 _031_
rlabel metal1 6302 13328 6302 13328 0 _032_
rlabel metal1 5750 13498 5750 13498 0 _033_
rlabel metal1 7866 13430 7866 13430 0 _034_
rlabel metal1 9844 13362 9844 13362 0 _035_
rlabel metal1 9522 13396 9522 13396 0 _036_
rlabel metal1 8878 12342 8878 12342 0 _037_
rlabel metal1 11270 13294 11270 13294 0 _038_
rlabel metal2 11362 13532 11362 13532 0 _039_
rlabel metal1 10902 13430 10902 13430 0 _040_
rlabel via1 10442 12954 10442 12954 0 _041_
rlabel metal1 10488 11186 10488 11186 0 _042_
rlabel metal1 10005 12342 10005 12342 0 _043_
rlabel metal1 11224 11866 11224 11866 0 _044_
rlabel metal1 10005 11254 10005 11254 0 _045_
rlabel metal1 6026 14484 6026 14484 0 _046_
rlabel metal1 9338 12750 9338 12750 0 bit_index\[0\]
rlabel metal2 7406 9690 7406 9690 0 bit_index\[1\]
rlabel metal1 6348 11662 6348 11662 0 bit_index\[2\]
rlabel metal2 6486 12563 6486 12563 0 clk
rlabel metal1 6601 12750 6601 12750 0 clknet_0_clk
rlabel metal1 4784 13906 4784 13906 0 clknet_1_0__leaf_clk
rlabel metal1 10994 14518 10994 14518 0 clknet_1_1__leaf_clk
rlabel metal2 8510 578 8510 578 0 comp
rlabel metal1 14812 11866 14812 11866 0 data_out[0]
rlabel metal1 12972 12954 12972 12954 0 data_out[1]
rlabel metal1 12650 14246 12650 14246 0 data_out[2]
rlabel metal1 10396 14042 10396 14042 0 data_out[3]
rlabel metal1 8694 15130 8694 15130 0 data_out[4]
rlabel metal2 7222 15140 7222 15140 0 data_out[5]
rlabel metal1 5934 14586 5934 14586 0 data_out[6]
rlabel metal1 4876 14586 4876 14586 0 data_out[7]
rlabel metal2 5566 13532 5566 13532 0 net1
rlabel metal1 8326 11254 8326 11254 0 net10
rlabel metal1 6486 11730 6486 11730 0 net11
rlabel metal2 4646 14620 4646 14620 0 net2
rlabel metal1 2714 12206 2714 12206 0 net3
rlabel metal2 7682 13532 7682 13532 0 net4
rlabel metal2 9982 11390 9982 11390 0 net5
rlabel metal1 7176 13838 7176 13838 0 net6
rlabel metal1 6532 12274 6532 12274 0 net7
rlabel metal1 6486 9520 6486 9520 0 net8
rlabel metal2 6302 10404 6302 10404 0 net9
rlabel metal2 12742 11492 12742 11492 0 out_data\[0\]
rlabel metal2 12742 12580 12742 12580 0 out_data\[1\]
rlabel metal1 12788 14450 12788 14450 0 out_data\[2\]
rlabel metal2 10534 14042 10534 14042 0 out_data\[3\]
rlabel metal2 8510 14076 8510 14076 0 out_data\[4\]
rlabel metal2 6394 14246 6394 14246 0 out_data\[5\]
rlabel metal1 7084 11662 7084 11662 0 out_data\[6\]
rlabel metal1 5934 13294 5934 13294 0 out_data\[7\]
rlabel metal2 1058 15317 1058 15317 0 reset
rlabel metal1 8464 12750 8464 12750 0 state
<< properties >>
string FIXED_BBOX 0 0 16000 16000
<< end >>
