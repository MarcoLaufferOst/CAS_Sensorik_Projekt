magic
tech sky130A
magscale 1 2
timestamp 1736799799
<< mvnmos >>
rect -629 -300 -29 300
rect 29 -300 629 300
<< mvndiff >>
rect -687 288 -629 300
rect -687 -288 -675 288
rect -641 -288 -629 288
rect -687 -300 -629 -288
rect -29 288 29 300
rect -29 -288 -17 288
rect 17 -288 29 288
rect -29 -300 29 -288
rect 629 288 687 300
rect 629 -288 641 288
rect 675 -288 687 288
rect 629 -300 687 -288
<< mvndiffc >>
rect -675 -288 -641 288
rect -17 -288 17 288
rect 641 -288 675 288
<< poly >>
rect -629 372 -29 388
rect -629 338 -613 372
rect -45 338 -29 372
rect -629 300 -29 338
rect 29 372 629 388
rect 29 338 45 372
rect 613 338 629 372
rect 29 300 629 338
rect -629 -338 -29 -300
rect -629 -372 -613 -338
rect -45 -372 -29 -338
rect -629 -388 -29 -372
rect 29 -338 629 -300
rect 29 -372 45 -338
rect 613 -372 629 -338
rect 29 -388 629 -372
<< polycont >>
rect -613 338 -45 372
rect 45 338 613 372
rect -613 -372 -45 -338
rect 45 -372 613 -338
<< locali >>
rect -629 338 -613 372
rect -45 338 -29 372
rect 29 338 45 372
rect 613 338 629 372
rect -675 288 -641 304
rect -675 -304 -641 -288
rect -17 288 17 304
rect -17 -304 17 -288
rect 641 288 675 304
rect 641 -304 675 -288
rect -629 -372 -613 -338
rect -45 -372 -29 -338
rect 29 -372 45 -338
rect 613 -372 629 -338
<< viali >>
rect -613 338 -45 372
rect 45 338 613 372
rect -675 -288 -641 288
rect -17 -288 17 288
rect 641 -288 675 288
rect -613 -372 -45 -338
rect 45 -372 613 -338
<< metal1 >>
rect -625 372 -33 378
rect -625 338 -613 372
rect -45 338 -33 372
rect -625 332 -33 338
rect 33 372 625 378
rect 33 338 45 372
rect 613 338 625 372
rect 33 332 625 338
rect -681 288 -635 300
rect -681 -288 -675 288
rect -641 -288 -635 288
rect -681 -300 -635 -288
rect -23 288 23 300
rect -23 -288 -17 288
rect 17 -288 23 288
rect -23 -300 23 -288
rect 635 288 681 300
rect 635 -288 641 288
rect 675 -288 681 288
rect 635 -300 681 -288
rect -625 -338 -33 -332
rect -625 -372 -613 -338
rect -45 -372 -33 -338
rect -625 -378 -33 -372
rect 33 -338 625 -332
rect 33 -372 45 -338
rect 613 -372 625 -338
rect 33 -378 625 -372
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 3.0 l 3.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
