magic
tech sky130A
magscale 1 2
timestamp 1736255080
<< nwell >>
rect 1880 1129 2790 2600
rect 1880 1124 2206 1129
rect 1880 975 2191 1124
rect 2320 1119 2790 1129
rect 2320 980 2510 1119
rect 2310 975 2510 980
rect 1880 970 2510 975
rect 2623 970 2790 1119
rect 1880 -610 2790 970
<< mvpsubdiff >>
rect 1300 2430 1790 2440
rect 1300 2390 1390 2430
rect 1700 2390 1790 2430
rect 1300 2380 1790 2390
rect 1300 2350 1360 2380
rect 1300 -460 1310 2350
rect 1350 -460 1360 2350
rect 1300 -490 1360 -460
rect 1730 2350 1790 2380
rect 1730 -460 1740 2350
rect 1780 -460 1790 2350
rect 1730 -490 1790 -460
rect 1300 -500 1790 -490
rect 1300 -540 1380 -500
rect 1710 -540 1790 -500
rect 1300 -550 1790 -540
<< mvnsubdiff >>
rect 1950 2420 2720 2430
rect 1950 2380 2040 2420
rect 2630 2380 2720 2420
rect 1950 2370 2720 2380
rect 1950 2340 2010 2370
rect 1950 -450 1960 2340
rect 2000 -450 2010 2340
rect 1950 -480 2010 -450
rect 2660 2340 2720 2370
rect 2660 -450 2670 2340
rect 2710 -450 2720 2340
rect 2660 -480 2720 -450
rect 1950 -490 2720 -480
rect 1950 -530 2040 -490
rect 2630 -530 2720 -490
rect 1950 -540 2720 -530
<< mvpsubdiffcont >>
rect 1390 2390 1700 2430
rect 1310 -460 1350 2350
rect 1740 -460 1780 2350
rect 1380 -540 1710 -500
<< mvnsubdiffcont >>
rect 2040 2380 2630 2420
rect 1960 -450 2000 2340
rect 2670 -450 2710 2340
rect 2040 -530 2630 -490
<< locali >>
rect 1310 2390 1390 2430
rect 1700 2390 1780 2430
rect 1310 2350 1350 2390
rect 1310 -500 1350 -460
rect 1740 2350 1780 2390
rect 1740 -500 1780 -460
rect 1310 -540 1380 -500
rect 1710 -540 1780 -500
rect 1960 2380 2040 2420
rect 2630 2380 2710 2420
rect 1960 2340 2000 2380
rect 1960 -490 2000 -450
rect 2670 2340 2710 2380
rect 2670 -490 2710 -450
rect 1960 -530 2040 -490
rect 2630 -530 2710 -490
<< viali >>
rect 1390 2390 1700 2430
rect 1310 -460 1350 2350
rect 1740 -460 1780 2350
rect 1380 -540 1710 -500
rect 2040 2380 2630 2420
rect 1960 -450 2000 2340
rect 2670 -450 2710 2340
rect 2040 -530 2630 -490
<< metal1 >>
rect 1200 2830 9610 2870
rect 1200 2670 2840 2830
rect 2940 2670 9610 2830
rect 1200 2470 9610 2670
rect 1300 2430 1790 2440
rect 1300 2390 1390 2430
rect 1700 2390 1790 2430
rect 1300 2380 1790 2390
rect 1300 2350 1360 2380
rect 1300 -460 1310 2350
rect 1350 -460 1360 2350
rect 1730 2350 1790 2380
rect 1588 990 1598 1190
rect 1656 990 1666 1190
rect 1430 790 1440 890
rect 1498 790 1508 890
rect 1488 217 1498 277
rect 1598 217 1608 277
rect 1488 -186 1498 -126
rect 1598 -186 1608 -126
rect 1430 -360 1440 -260
rect 1498 -360 1508 -260
rect 1300 -490 1360 -460
rect 1419 -490 1519 -396
rect 1588 -410 1598 -310
rect 1656 -410 1666 -310
rect 1730 -460 1740 2350
rect 1780 -460 1790 2350
rect 1730 -490 1790 -460
rect 1300 -500 1790 -490
rect 1300 -540 1380 -500
rect 1710 -540 1790 -500
rect 1950 2420 2720 2470
rect 1950 2380 2040 2420
rect 2630 2380 2720 2420
rect 1950 2370 2720 2380
rect 1950 2340 2010 2370
rect 1950 -450 1960 2340
rect 2000 -450 2010 2340
rect 2660 2340 2720 2370
rect 2214 990 2224 1190
rect 2283 990 2293 1190
rect 2530 990 2540 1190
rect 2598 990 2608 1190
rect 2056 790 2066 890
rect 2124 790 2134 890
rect 2372 790 2382 890
rect 2440 790 2450 890
rect 2114 220 2124 280
rect 2224 220 2234 280
rect 2272 220 2282 280
rect 2382 220 2392 280
rect 2430 220 2440 280
rect 2540 220 2550 280
rect 2114 -190 2124 -130
rect 2224 -190 2234 -130
rect 2272 -190 2282 -130
rect 2382 -190 2392 -130
rect 2430 -190 2440 -130
rect 2540 -190 2550 -130
rect 2056 -410 2066 -310
rect 2124 -410 2134 -310
rect 2214 -424 2224 -324
rect 2282 -424 2292 -324
rect 2372 -424 2382 -324
rect 2440 -424 2450 -324
rect 2530 -424 2540 -324
rect 2598 -424 2608 -324
rect 1950 -480 2010 -450
rect 2660 -450 2670 2340
rect 2710 -450 2720 2340
rect 2660 -480 2720 -450
rect 1950 -490 2720 -480
rect 1950 -530 2040 -490
rect 2630 -530 2720 -490
rect 1950 -540 2720 -530
rect 1300 -570 1790 -540
rect 1200 -690 9610 -570
rect 1200 -850 1419 -690
rect 1519 -700 9610 -690
rect 1519 -850 2640 -700
rect 1200 -900 2640 -850
rect 2840 -900 9610 -700
rect 1200 -970 9610 -900
<< via1 >>
rect 2840 2670 2940 2830
rect 1598 990 1656 1190
rect 1440 790 1498 890
rect 1498 217 1598 277
rect 1498 -186 1598 -126
rect 1440 -360 1498 -260
rect 1598 -410 1656 -310
rect 2224 990 2283 1190
rect 2540 990 2598 1190
rect 2066 790 2124 890
rect 2382 790 2440 890
rect 2124 220 2224 280
rect 2282 220 2382 280
rect 2440 220 2540 280
rect 2124 -190 2224 -130
rect 2282 -190 2382 -130
rect 2440 -190 2540 -130
rect 2066 -410 2124 -310
rect 2224 -424 2282 -324
rect 2382 -424 2440 -324
rect 2540 -424 2598 -324
rect 1419 -850 1519 -690
rect 2640 -900 2840 -700
<< metal2 >>
rect 2840 2830 2940 2840
rect 1598 1190 1656 1200
rect 1598 980 1656 990
rect 2224 1190 2283 1200
rect 2224 980 2283 990
rect 2540 1190 2598 1200
rect 2540 980 2598 990
rect 1440 890 1498 900
rect 1440 780 1498 790
rect 2066 890 2124 900
rect 2066 780 2124 790
rect 2382 890 2440 900
rect 2382 780 2440 790
rect 2640 300 2740 310
rect 1498 277 1598 287
rect 1498 100 1598 217
rect 2124 280 2224 290
rect 2124 210 2224 220
rect 2282 280 2382 290
rect 2282 210 2382 220
rect 2440 280 2540 290
rect 2440 210 2540 220
rect 1498 -10 1598 0
rect 1790 100 1890 110
rect 1790 -110 1890 0
rect 1498 -126 1598 -116
rect 1498 -196 1598 -186
rect 2124 -130 2224 -120
rect 2124 -200 2224 -190
rect 2282 -130 2382 -120
rect 2282 -200 2382 -190
rect 2440 -130 2540 -120
rect 2440 -200 2540 -190
rect 1790 -220 1890 -210
rect 1440 -260 1498 -250
rect 1419 -360 1440 -260
rect 1498 -360 1519 -260
rect 1419 -690 1519 -360
rect 1598 -310 1656 -300
rect 1598 -420 1656 -410
rect 2066 -310 2124 -300
rect 2640 -310 2740 200
rect 2224 -324 2282 -314
rect 2382 -324 2440 -314
rect 2066 -420 2124 -410
rect 2203 -424 2224 -324
rect 2282 -424 2303 -324
rect 2203 -510 2303 -424
rect 2382 -434 2440 -424
rect 2510 -324 2610 -310
rect 2510 -424 2540 -324
rect 2598 -424 2610 -324
rect 2640 -420 2740 -410
rect 2203 -620 2303 -610
rect 2510 -510 2610 -424
rect 2510 -620 2610 -610
rect 2840 -510 2940 2670
rect 2840 -620 2940 -610
rect 1419 -860 1519 -850
rect 2640 -700 2840 -690
rect 2640 -910 2840 -900
<< via2 >>
rect 1598 990 1656 1190
rect 2224 990 2283 1190
rect 2540 990 2598 1190
rect 1440 790 1498 890
rect 2066 790 2124 890
rect 2382 790 2440 890
rect 2124 220 2224 280
rect 2282 220 2382 280
rect 2440 220 2540 280
rect 2640 200 2740 300
rect 1498 0 1598 100
rect 1790 0 1890 100
rect 1498 -186 1598 -126
rect 1790 -210 1890 -110
rect 2124 -190 2224 -130
rect 2282 -190 2382 -130
rect 2440 -190 2540 -130
rect 1598 -410 1656 -310
rect 2066 -410 2124 -310
rect 2382 -424 2440 -324
rect 2640 -410 2740 -310
rect 2203 -610 2303 -510
rect 2510 -610 2610 -510
rect 2840 -610 2940 -510
rect 2640 -900 2840 -700
<< metal3 >>
rect 1588 1190 1666 1195
rect 2214 1190 2293 1195
rect 2530 1190 2608 1195
rect 1420 990 1598 1190
rect 1656 990 2224 1190
rect 2283 990 2540 1190
rect 2598 990 2840 1190
rect 2940 990 2950 1190
rect 9190 990 9200 1190
rect 9400 990 9610 1190
rect 1588 985 1666 990
rect 2214 985 2293 990
rect 2530 985 2608 990
rect 1430 890 1508 895
rect 2056 890 2134 895
rect 2372 890 2450 895
rect 1200 790 1440 890
rect 1498 790 2066 890
rect 2124 790 2382 890
rect 2440 790 2610 890
rect 1430 785 1508 790
rect 2056 785 2134 790
rect 2372 785 2450 790
rect 2630 300 2750 305
rect 1300 280 2640 300
rect 1300 220 2124 280
rect 2224 220 2282 280
rect 2382 220 2440 280
rect 2540 220 2640 280
rect 1300 200 2640 220
rect 2740 200 2750 300
rect 2630 195 2750 200
rect 1488 100 1608 105
rect 1780 100 1900 105
rect 1200 0 1498 100
rect 1598 0 1790 100
rect 1890 0 2640 100
rect 1488 -5 1608 0
rect 1780 -5 1900 0
rect 1780 -110 1900 -105
rect 1300 -126 1790 -110
rect 1300 -186 1498 -126
rect 1598 -186 1790 -126
rect 1300 -210 1790 -186
rect 1890 -130 2640 -110
rect 1890 -190 2124 -130
rect 2224 -190 2282 -130
rect 2382 -190 2440 -130
rect 2540 -190 2640 -130
rect 1890 -210 2640 -190
rect 1780 -215 1900 -210
rect 1588 -310 1666 -305
rect 2056 -310 2134 -305
rect 2630 -310 2750 -305
rect 1580 -410 1598 -310
rect 1656 -410 2066 -310
rect 2124 -324 2640 -310
rect 2124 -410 2382 -324
rect 1588 -415 1666 -410
rect 2056 -415 2134 -410
rect 2372 -424 2382 -410
rect 2440 -410 2640 -324
rect 2740 -410 2790 -310
rect 2440 -424 2450 -410
rect 2630 -415 2750 -410
rect 2372 -429 2450 -424
rect 2193 -510 2313 -505
rect 2500 -510 2620 -505
rect 2830 -510 2950 -505
rect 2160 -610 2203 -510
rect 2303 -610 2510 -510
rect 2610 -610 2840 -510
rect 2940 -610 2950 -510
rect 2193 -615 2313 -610
rect 2500 -615 2620 -610
rect 2830 -615 2950 -610
rect 2630 -700 2850 -695
rect 2630 -900 2640 -700
rect 2840 -900 3560 -700
rect 2630 -905 2850 -900
<< via3 >>
rect 2840 990 2940 1190
rect 9200 990 9400 1190
<< metal4 >>
rect 2839 1190 2941 1191
rect 9199 1190 9401 1191
rect 2839 990 2840 1190
rect 2940 990 9200 1190
rect 9400 990 9401 1190
rect 2839 989 2941 990
rect 9199 989 9401 990
use sky130_fd_pr__cap_mim_m3_1_9ZMSDV  XC1
timestamp 1736253881
transform 0 1 6070 1 0 916
box -1886 -3040 1886 3040
use sky130_fd_pr__nfet_g5v0d10v5_SMV9TY  XM3
timestamp 1736238736
transform 1 0 1548 0 1 -283
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_PEM9WF  XM4
timestamp 1736238736
transform -1 0 2332 0 1 -288
box -332 -202 332 164
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM5
timestamp 1736238736
transform -1 0 1548 0 -1 1274
box -108 -1057 108 1057
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM6
timestamp 1736238736
transform -1 0 2332 0 -1 1278
box -332 -1102 332 1064
<< labels >>
flabel metal1 1200 -970 1300 -870 0 FreeSans 160 0 0 0 vssa
port 6 nsew
flabel metal3 1200 0 1300 100 0 FreeSans 160 0 0 0 sample
port 1 nsew
flabel metal1 1200 2770 1300 2870 0 FreeSans 160 0 0 0 vdda
port 5 nsew
flabel metal3 1200 790 1300 890 0 FreeSans 160 0 0 0 vin
port 18 nsew
flabel metal3 9510 990 9610 1090 0 FreeSans 160 0 0 0 vout
port 17 nsew
<< end >>
