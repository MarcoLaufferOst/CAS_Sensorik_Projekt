magic
tech sky130A
magscale 1 2
timestamp 1736799598
<< error_p >>
rect -753 -166 -723 166
rect -687 -100 -657 100
rect 657 -100 687 100
rect 723 -166 753 166
<< nwell >>
rect -723 -200 723 200
<< mvpmos >>
rect -629 -100 -29 100
rect 29 -100 629 100
<< mvpdiff >>
rect -687 88 -629 100
rect -687 -88 -675 88
rect -641 -88 -629 88
rect -687 -100 -629 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 629 88 687 100
rect 629 -88 641 88
rect 675 -88 687 88
rect 629 -100 687 -88
<< mvpdiffc >>
rect -675 -88 -641 88
rect -17 -88 17 88
rect 641 -88 675 88
<< poly >>
rect -629 181 -29 197
rect -629 147 -613 181
rect -45 147 -29 181
rect -629 100 -29 147
rect 29 181 629 197
rect 29 147 45 181
rect 613 147 629 181
rect 29 100 629 147
rect -629 -147 -29 -100
rect -629 -181 -613 -147
rect -45 -181 -29 -147
rect -629 -197 -29 -181
rect 29 -147 629 -100
rect 29 -181 45 -147
rect 613 -181 629 -147
rect 29 -197 629 -181
<< polycont >>
rect -613 147 -45 181
rect 45 147 613 181
rect -613 -181 -45 -147
rect 45 -181 613 -147
<< locali >>
rect -629 147 -613 181
rect -45 147 -29 181
rect 29 147 45 181
rect 613 147 629 181
rect -675 88 -641 104
rect -675 -104 -641 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 641 88 675 104
rect 641 -104 675 -88
rect -629 -181 -613 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 613 -181 629 -147
<< viali >>
rect -613 147 -45 181
rect 45 147 613 181
rect -675 -88 -641 88
rect -17 -88 17 88
rect 641 -88 675 88
rect -613 -181 -45 -147
rect 45 -181 613 -147
<< metal1 >>
rect -625 181 -33 187
rect -625 147 -613 181
rect -45 147 -33 181
rect -625 141 -33 147
rect 33 181 625 187
rect 33 147 45 181
rect 613 147 625 181
rect 33 141 625 147
rect -681 88 -635 100
rect -681 -88 -675 88
rect -641 -88 -635 88
rect -681 -100 -635 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 635 88 681 100
rect 635 -88 641 88
rect 675 -88 681 88
rect 635 -100 681 -88
rect -625 -147 -33 -141
rect -625 -181 -613 -147
rect -45 -181 -33 -147
rect -625 -187 -33 -181
rect 33 -147 625 -141
rect 33 -181 45 -147
rect 613 -181 625 -147
rect 33 -187 625 -181
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 1 l 3.0 m 1 nf 2 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
