magic
tech sky130A
magscale 1 2
timestamp 1735905635
<< mvnmos >>
rect -487 -1750 -287 1750
rect -229 -1750 -29 1750
rect 29 -1750 229 1750
rect 287 -1750 487 1750
<< mvndiff >>
rect -545 1738 -487 1750
rect -545 -1738 -533 1738
rect -499 -1738 -487 1738
rect -545 -1750 -487 -1738
rect -287 1738 -229 1750
rect -287 -1738 -275 1738
rect -241 -1738 -229 1738
rect -287 -1750 -229 -1738
rect -29 1738 29 1750
rect -29 -1738 -17 1738
rect 17 -1738 29 1738
rect -29 -1750 29 -1738
rect 229 1738 287 1750
rect 229 -1738 241 1738
rect 275 -1738 287 1738
rect 229 -1750 287 -1738
rect 487 1738 545 1750
rect 487 -1738 499 1738
rect 533 -1738 545 1738
rect 487 -1750 545 -1738
<< mvndiffc >>
rect -533 -1738 -499 1738
rect -275 -1738 -241 1738
rect -17 -1738 17 1738
rect 241 -1738 275 1738
rect 499 -1738 533 1738
<< poly >>
rect -487 1822 -287 1838
rect -487 1788 -471 1822
rect -303 1788 -287 1822
rect -487 1750 -287 1788
rect -229 1822 -29 1838
rect -229 1788 -213 1822
rect -45 1788 -29 1822
rect -229 1750 -29 1788
rect 29 1822 229 1838
rect 29 1788 45 1822
rect 213 1788 229 1822
rect 29 1750 229 1788
rect 287 1822 487 1838
rect 287 1788 303 1822
rect 471 1788 487 1822
rect 287 1750 487 1788
rect -487 -1788 -287 -1750
rect -487 -1822 -471 -1788
rect -303 -1822 -287 -1788
rect -487 -1838 -287 -1822
rect -229 -1788 -29 -1750
rect -229 -1822 -213 -1788
rect -45 -1822 -29 -1788
rect -229 -1838 -29 -1822
rect 29 -1788 229 -1750
rect 29 -1822 45 -1788
rect 213 -1822 229 -1788
rect 29 -1838 229 -1822
rect 287 -1788 487 -1750
rect 287 -1822 303 -1788
rect 471 -1822 487 -1788
rect 287 -1838 487 -1822
<< polycont >>
rect -471 1788 -303 1822
rect -213 1788 -45 1822
rect 45 1788 213 1822
rect 303 1788 471 1822
rect -471 -1822 -303 -1788
rect -213 -1822 -45 -1788
rect 45 -1822 213 -1788
rect 303 -1822 471 -1788
<< locali >>
rect -487 1788 -471 1822
rect -303 1788 -287 1822
rect -229 1788 -213 1822
rect -45 1788 -29 1822
rect 29 1788 45 1822
rect 213 1788 229 1822
rect 287 1788 303 1822
rect 471 1788 487 1822
rect -533 1738 -499 1754
rect -533 -1754 -499 -1738
rect -275 1738 -241 1754
rect -275 -1754 -241 -1738
rect -17 1738 17 1754
rect -17 -1754 17 -1738
rect 241 1738 275 1754
rect 241 -1754 275 -1738
rect 499 1738 533 1754
rect 499 -1754 533 -1738
rect -487 -1822 -471 -1788
rect -303 -1822 -287 -1788
rect -229 -1822 -213 -1788
rect -45 -1822 -29 -1788
rect 29 -1822 45 -1788
rect 213 -1822 229 -1788
rect 287 -1822 303 -1788
rect 471 -1822 487 -1788
<< viali >>
rect -471 1788 -303 1822
rect -213 1788 -45 1822
rect 45 1788 213 1822
rect 303 1788 471 1822
rect -533 -1738 -499 1738
rect -275 -1738 -241 1738
rect -17 -1738 17 1738
rect 241 -1738 275 1738
rect 499 -1738 533 1738
rect -471 -1822 -303 -1788
rect -213 -1822 -45 -1788
rect 45 -1822 213 -1788
rect 303 -1822 471 -1788
<< metal1 >>
rect -483 1822 -291 1828
rect -483 1788 -471 1822
rect -303 1788 -291 1822
rect -483 1782 -291 1788
rect -225 1822 -33 1828
rect -225 1788 -213 1822
rect -45 1788 -33 1822
rect -225 1782 -33 1788
rect 33 1822 225 1828
rect 33 1788 45 1822
rect 213 1788 225 1822
rect 33 1782 225 1788
rect 291 1822 483 1828
rect 291 1788 303 1822
rect 471 1788 483 1822
rect 291 1782 483 1788
rect -539 1738 -493 1750
rect -539 -1738 -533 1738
rect -499 -1738 -493 1738
rect -539 -1750 -493 -1738
rect -281 1738 -235 1750
rect -281 -1738 -275 1738
rect -241 -1738 -235 1738
rect -281 -1750 -235 -1738
rect -23 1738 23 1750
rect -23 -1738 -17 1738
rect 17 -1738 23 1738
rect -23 -1750 23 -1738
rect 235 1738 281 1750
rect 235 -1738 241 1738
rect 275 -1738 281 1738
rect 235 -1750 281 -1738
rect 493 1738 539 1750
rect 493 -1738 499 1738
rect 533 -1738 539 1738
rect 493 -1750 539 -1738
rect -483 -1788 -291 -1782
rect -483 -1822 -471 -1788
rect -303 -1822 -291 -1788
rect -483 -1828 -291 -1822
rect -225 -1788 -33 -1782
rect -225 -1822 -213 -1788
rect -45 -1822 -33 -1788
rect -225 -1828 -33 -1822
rect 33 -1788 225 -1782
rect 33 -1822 45 -1788
rect 213 -1822 225 -1788
rect 33 -1828 225 -1822
rect 291 -1788 483 -1782
rect 291 -1822 303 -1788
rect 471 -1822 483 -1788
rect 291 -1828 483 -1822
<< properties >>
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 17.5 l 1.0 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
