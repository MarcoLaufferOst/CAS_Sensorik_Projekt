magic
tech sky130A
magscale 1 2
timestamp 1736447341
<< nwell >>
rect 1530 -5400 6190 -3890
rect 1530 -7220 6190 -6350
rect 1530 -7710 3910 -7220
rect 3960 -7710 6190 -7220
rect 1530 -7860 6190 -7710
rect 1550 -8970 6190 -8810
rect 1550 -9030 1790 -8970
rect 1550 -9500 1740 -9030
rect 1800 -9500 6190 -8970
rect 1550 -9720 6190 -9500
rect 4100 -9900 6190 -9720
rect 4100 -9960 4410 -9900
rect 4560 -9910 4680 -9900
rect 4830 -9960 6190 -9900
rect 4100 -10470 6190 -9960
<< mvpsubdiff >>
rect 1600 -3320 6120 -3310
rect 1600 -3360 1670 -3320
rect 6050 -3360 6120 -3320
rect 1600 -3370 6120 -3360
rect 1600 -3740 1660 -3370
rect 6060 -3740 6120 -3370
rect 1600 -3750 6120 -3740
rect 1600 -3790 1670 -3750
rect 6050 -3790 6120 -3750
rect 1600 -3800 6120 -3790
rect 1600 -5500 6120 -5490
rect 1600 -5540 1670 -5500
rect 6050 -5540 6120 -5500
rect 1600 -5550 6120 -5540
rect 1600 -5560 1680 -5550
rect 1600 -6200 1660 -5560
rect 6060 -6200 6120 -5550
rect 1600 -6210 6120 -6200
rect 1600 -6250 1670 -6210
rect 6050 -6250 6120 -6210
rect 1600 -6260 6120 -6250
rect 1600 -7960 2710 -7950
rect 2960 -7960 6120 -7950
rect 1600 -8000 1670 -7960
rect 6050 -8000 6120 -7960
rect 1600 -8010 6120 -8000
rect 1600 -8660 1660 -8010
rect 6060 -8660 6120 -8010
rect 1600 -8670 6120 -8660
rect 1600 -8710 1670 -8670
rect 6050 -8710 6120 -8670
rect 1600 -8720 6120 -8710
rect 1620 -9820 4010 -9810
rect 1620 -9860 1670 -9820
rect 3960 -9860 4010 -9820
rect 1620 -9870 4010 -9860
rect 1620 -10340 1680 -9870
rect 3950 -10340 4010 -9870
rect 1620 -10350 4010 -10340
rect 1620 -10390 1670 -10350
rect 3960 -10390 4010 -10350
rect 1620 -10400 4010 -10390
<< mvnsubdiff >>
rect 1600 -3970 6120 -3960
rect 1600 -4010 1670 -3970
rect 6050 -4010 6120 -3970
rect 1600 -4020 6120 -4010
rect 1600 -5270 1660 -4020
rect 6060 -5270 6120 -4020
rect 1600 -5280 6120 -5270
rect 1600 -5320 1670 -5280
rect 6050 -5320 6120 -5280
rect 1600 -5330 6120 -5320
rect 1600 -6430 6120 -6420
rect 1600 -6470 1670 -6430
rect 6050 -6470 6120 -6430
rect 1600 -6480 6120 -6470
rect 1600 -7730 1660 -6480
rect 6060 -7730 6120 -6480
rect 1600 -7740 6120 -7730
rect 1600 -7780 1670 -7740
rect 6050 -7780 6120 -7740
rect 1600 -7790 6120 -7780
rect 1620 -8890 6120 -8880
rect 1620 -8930 1670 -8890
rect 6050 -8930 6120 -8890
rect 1620 -8940 6120 -8930
rect 1620 -9590 1680 -8940
rect 1620 -9600 4230 -9590
rect 1620 -9640 1670 -9600
rect 4180 -9640 4230 -9600
rect 1620 -9650 4230 -9640
rect 4170 -10340 4230 -9650
rect 6060 -10340 6120 -8940
rect 4170 -10350 6120 -10340
rect 4170 -10390 4220 -10350
rect 6050 -10390 6120 -10350
rect 4170 -10400 6120 -10390
<< mvpsubdiffcont >>
rect 1670 -3360 6050 -3320
rect 1670 -3790 6050 -3750
rect 1670 -5540 6050 -5500
rect 1670 -6250 6050 -6210
rect 1670 -8000 6050 -7960
rect 1670 -8710 6050 -8670
rect 1670 -9860 3960 -9820
rect 1670 -10390 3960 -10350
<< mvnsubdiffcont >>
rect 1670 -4010 6050 -3970
rect 1670 -5320 6050 -5280
rect 1670 -6470 6050 -6430
rect 1670 -7780 6050 -7740
rect 1670 -8930 6050 -8890
rect 1670 -9640 4180 -9600
rect 4220 -10390 6050 -10350
<< locali >>
rect 1610 -3360 1670 -3320
rect 6050 -3360 6110 -3320
rect 1610 -3750 1650 -3360
rect 6070 -3750 6110 -3360
rect 1610 -3790 1670 -3750
rect 6050 -3790 6110 -3750
rect 1610 -4010 1670 -3970
rect 6050 -4010 6110 -3970
rect 1610 -5280 1650 -4010
rect 6070 -5280 6110 -4010
rect 1610 -5320 1670 -5280
rect 6050 -5320 6110 -5280
rect 1610 -5550 1670 -5500
rect 6050 -5540 6110 -5500
rect 1610 -6200 1650 -5550
rect 1610 -6250 1670 -6200
rect 6070 -6210 6110 -5540
rect 6050 -6250 6110 -6210
rect 1610 -6470 1670 -6430
rect 6050 -6470 6110 -6430
rect 1610 -7740 1650 -6470
rect 6070 -7740 6110 -6470
rect 1610 -7780 1670 -7740
rect 6050 -7780 6110 -7740
rect 1610 -8000 1670 -7960
rect 6050 -8000 6110 -7960
rect 1610 -8670 1650 -8000
rect 6070 -8670 6110 -8000
rect 1610 -8710 1670 -8670
rect 6050 -8710 6110 -8670
rect 1630 -9640 1670 -8890
rect 6050 -8930 6110 -8890
rect 1630 -10390 1670 -9820
rect 3960 -10390 4000 -9820
rect 4180 -10390 4220 -9600
rect 6070 -10350 6110 -8930
rect 6050 -10390 6110 -10350
<< viali >>
rect 1670 -3360 6050 -3320
rect 1670 -3790 6050 -3750
rect 1670 -4010 6050 -3970
rect 1670 -5320 6050 -5280
rect 1670 -5540 6050 -5500
rect 1670 -6250 6050 -6210
rect 1670 -6470 6050 -6430
rect 1670 -7780 6050 -7740
rect 1670 -8000 6050 -7960
rect 1670 -8710 6050 -8670
rect 1670 -8930 6050 -8890
rect 1670 -9640 4180 -9600
rect 1670 -9860 3960 -9820
rect 1670 -10390 3960 -10350
rect 4220 -10390 6050 -10350
<< metal1 >>
rect 1150 -3320 6130 -3170
rect 1150 -3360 1670 -3320
rect 6050 -3360 6130 -3320
rect 1150 -3370 6130 -3360
rect 1150 -5360 1550 -3370
rect 1600 -3740 1660 -3370
rect 1810 -3490 5910 -3400
rect 1690 -3600 1700 -3500
rect 1770 -3600 1780 -3500
rect 5940 -3600 5950 -3500
rect 6020 -3600 6030 -3500
rect 2350 -3660 2360 -3600
rect 2460 -3660 2470 -3600
rect 5210 -3660 5220 -3600
rect 5320 -3660 5330 -3600
rect 6060 -3740 6120 -3370
rect 1600 -3750 6120 -3740
rect 1600 -3790 1670 -3750
rect 6050 -3790 6120 -3750
rect 1600 -3800 6120 -3790
rect 6160 -3830 6560 -3170
rect 1590 -3970 6560 -3830
rect 1590 -4010 1670 -3970
rect 6050 -4010 6560 -3970
rect 1590 -4030 6560 -4010
rect 1600 -5270 1660 -4030
rect 2350 -4140 2360 -4080
rect 2460 -4140 2470 -4080
rect 5210 -4140 5220 -4080
rect 5320 -4140 5330 -4080
rect 1690 -4300 1760 -4140
rect 2950 -4300 2960 -4240
rect 3060 -4300 3070 -4240
rect 4450 -4300 4460 -4240
rect 4560 -4300 4570 -4240
rect 5960 -4300 6030 -4140
rect 1690 -4400 1700 -4300
rect 1770 -4400 1780 -4300
rect 5950 -4400 5960 -4300
rect 6020 -4400 6030 -4300
rect 1690 -4560 1760 -4400
rect 2350 -4460 2360 -4400
rect 2460 -4460 2470 -4400
rect 5210 -4460 5220 -4400
rect 5320 -4460 5330 -4400
rect 5960 -4560 6030 -4400
rect 2950 -4620 2960 -4560
rect 3060 -4620 3070 -4560
rect 4450 -4620 4460 -4560
rect 4560 -4620 4570 -4560
rect 2950 -4740 2960 -4680
rect 3060 -4740 3070 -4680
rect 4450 -4740 4460 -4680
rect 4560 -4740 4570 -4680
rect 1690 -4900 1760 -4740
rect 2350 -4900 2360 -4840
rect 2460 -4900 2470 -4840
rect 5210 -4900 5220 -4840
rect 5320 -4900 5330 -4840
rect 5960 -4900 6030 -4750
rect 1690 -5000 1700 -4900
rect 1770 -5000 1780 -4900
rect 5950 -5000 5960 -4900
rect 6020 -5000 6030 -4900
rect 1690 -5160 1760 -5000
rect 2950 -5060 2960 -5000
rect 3060 -5060 3070 -5000
rect 4450 -5060 4460 -5000
rect 4560 -5060 4570 -5000
rect 5960 -5150 6030 -5000
rect 2350 -5220 2360 -5160
rect 2460 -5220 2470 -5160
rect 5210 -5220 5220 -5160
rect 5320 -5220 5330 -5160
rect 6060 -5270 6120 -4030
rect 1600 -5280 6120 -5270
rect 1600 -5320 1670 -5280
rect 6050 -5320 6120 -5280
rect 1600 -5330 6120 -5320
rect 1150 -5500 6130 -5360
rect 1150 -5540 1670 -5500
rect 6050 -5540 6130 -5500
rect 1150 -5560 6130 -5540
rect 1150 -7820 1550 -5560
rect 1600 -6200 1660 -5560
rect 2350 -5680 2360 -5620
rect 2460 -5680 2470 -5620
rect 5210 -5680 5220 -5620
rect 5320 -5680 5330 -5620
rect 1690 -5780 1700 -5680
rect 1770 -5780 1780 -5680
rect 5940 -5780 5950 -5680
rect 6020 -5780 6030 -5680
rect 1810 -5850 5900 -5790
rect 1810 -5950 5900 -5890
rect 1690 -6060 1700 -5960
rect 1770 -6060 1780 -5960
rect 5940 -6060 5950 -5960
rect 6020 -6060 6030 -5960
rect 2350 -6120 2360 -6060
rect 2460 -6120 2470 -6060
rect 5210 -6120 5220 -6060
rect 5320 -6120 5330 -6060
rect 6060 -6200 6120 -5560
rect 1600 -6210 6120 -6200
rect 1600 -6250 1670 -6210
rect 6050 -6250 6120 -6210
rect 1600 -6260 6120 -6250
rect 6160 -6290 6560 -4030
rect 1590 -6430 6560 -6290
rect 1590 -6470 1670 -6430
rect 6050 -6470 6560 -6430
rect 1590 -6490 6560 -6470
rect 1600 -7730 1660 -6490
rect 2350 -6600 2360 -6540
rect 2460 -6600 2470 -6540
rect 5210 -6600 5220 -6540
rect 5320 -6600 5330 -6540
rect 1690 -6760 1760 -6600
rect 2950 -6760 2960 -6700
rect 3060 -6760 3070 -6700
rect 4450 -6760 4460 -6700
rect 4560 -6760 4570 -6700
rect 5960 -6760 6030 -6600
rect 1690 -6860 1700 -6760
rect 1770 -6860 1780 -6760
rect 5950 -6860 5960 -6760
rect 6020 -6860 6030 -6760
rect 1690 -7020 1760 -6860
rect 2350 -6920 2360 -6860
rect 2460 -6920 2470 -6860
rect 5210 -6920 5220 -6860
rect 5320 -6920 5330 -6860
rect 5960 -7020 6030 -6860
rect 2950 -7080 2960 -7020
rect 3060 -7080 3070 -7020
rect 4450 -7080 4460 -7020
rect 4560 -7080 4570 -7020
rect 2950 -7200 2960 -7140
rect 3060 -7200 3070 -7140
rect 4450 -7200 4460 -7140
rect 4560 -7200 4570 -7140
rect 1690 -7360 1760 -7200
rect 2280 -7360 2290 -7300
rect 2390 -7360 2400 -7300
rect 5210 -7360 5220 -7300
rect 5320 -7360 5330 -7300
rect 5960 -7360 6030 -7210
rect 1690 -7460 1700 -7360
rect 1770 -7460 1780 -7360
rect 5950 -7460 5960 -7360
rect 6020 -7460 6030 -7360
rect 1690 -7620 1760 -7460
rect 2950 -7520 2960 -7460
rect 3060 -7520 3070 -7460
rect 4450 -7520 4460 -7460
rect 4560 -7520 4570 -7460
rect 5960 -7620 6030 -7460
rect 2280 -7680 2290 -7620
rect 2390 -7680 2400 -7620
rect 5210 -7680 5220 -7620
rect 5320 -7680 5330 -7620
rect 6060 -7730 6120 -6490
rect 1600 -7740 6120 -7730
rect 1600 -7780 1670 -7740
rect 6050 -7780 6120 -7740
rect 1600 -7790 6120 -7780
rect 1150 -7860 6130 -7820
rect 1150 -7880 2490 -7860
rect 1150 -7960 1890 -7880
rect 1990 -7960 2490 -7880
rect 2590 -7960 3090 -7860
rect 3190 -7960 6130 -7860
rect 1150 -8000 1670 -7960
rect 6050 -8000 6130 -7960
rect 1150 -8020 6130 -8000
rect 1150 -10430 1550 -8020
rect 1600 -8660 1660 -8020
rect 2280 -8140 2290 -8080
rect 2390 -8140 2400 -8080
rect 5210 -8140 5220 -8080
rect 5320 -8140 5330 -8080
rect 1690 -8240 1700 -8140
rect 1770 -8240 1780 -8140
rect 5940 -8240 5950 -8140
rect 6020 -8240 6030 -8140
rect 1810 -8300 5900 -8240
rect 3080 -8360 3800 -8330
rect 1880 -8420 1890 -8360
rect 1990 -8420 2000 -8360
rect 2480 -8420 2490 -8360
rect 2590 -8420 2600 -8360
rect 3080 -8420 3090 -8360
rect 3190 -8390 3800 -8360
rect 3190 -8420 3200 -8390
rect 5210 -8420 5220 -8360
rect 5320 -8420 5330 -8360
rect 1710 -8520 1720 -8420
rect 1790 -8520 1800 -8420
rect 2280 -8510 2290 -8420
rect 2350 -8510 2360 -8420
rect 2890 -8520 2900 -8420
rect 2960 -8520 2970 -8420
rect 3490 -8520 3500 -8420
rect 3560 -8520 3570 -8420
rect 5940 -8520 5950 -8420
rect 6020 -8520 6030 -8420
rect 1880 -8580 1890 -8520
rect 1990 -8580 2000 -8520
rect 2480 -8580 2490 -8520
rect 2590 -8580 2600 -8520
rect 3080 -8580 3090 -8520
rect 3190 -8580 3200 -8520
rect 3680 -8580 3690 -8520
rect 3790 -8580 3800 -8520
rect 5410 -8580 5420 -8520
rect 5520 -8580 5530 -8520
rect 6060 -8660 6120 -8020
rect 1600 -8670 6120 -8660
rect 1600 -8710 1670 -8670
rect 6050 -8710 6120 -8670
rect 1600 -8720 6120 -8710
rect 6160 -8750 6560 -6490
rect 1590 -8850 2090 -8750
rect 2190 -8770 6560 -8750
rect 2190 -8850 2690 -8770
rect 1590 -8870 2690 -8850
rect 2790 -8780 6560 -8770
rect 2790 -8870 3290 -8780
rect 1590 -8880 3290 -8870
rect 3390 -8800 6560 -8780
rect 3390 -8880 5020 -8800
rect 1590 -8890 5020 -8880
rect 5120 -8890 6560 -8800
rect 1590 -8930 1670 -8890
rect 6050 -8930 6560 -8890
rect 1590 -8950 6560 -8930
rect 1620 -9590 1680 -8950
rect 1720 -9160 1730 -9050
rect 1790 -9160 1800 -9050
rect 1880 -9060 1890 -9002
rect 1990 -9060 2000 -9002
rect 2480 -9060 2490 -9000
rect 2590 -9060 2600 -9000
rect 3080 -9060 3090 -9000
rect 3190 -9060 3200 -9000
rect 3680 -9060 3690 -9000
rect 3790 -9060 3800 -9000
rect 5210 -9060 5220 -9000
rect 5320 -9060 5330 -9000
rect 2290 -9150 2300 -9060
rect 2360 -9150 2370 -9060
rect 2900 -9160 2910 -9060
rect 2970 -9160 2980 -9060
rect 3490 -9160 3500 -9060
rect 3560 -9160 3570 -9060
rect 1720 -9320 1730 -9210
rect 1790 -9320 1800 -9210
rect 1840 -9220 2090 -9160
rect 2190 -9220 2200 -9160
rect 2400 -9220 2690 -9160
rect 2790 -9220 2800 -9160
rect 3010 -9220 3290 -9160
rect 3390 -9220 3400 -9160
rect 3600 -9220 3880 -9160
rect 5410 -9220 5420 -9160
rect 5520 -9220 5530 -9160
rect 5960 -9220 6030 -9070
rect 2290 -9310 2300 -9220
rect 2360 -9310 2370 -9220
rect 1720 -9480 1730 -9370
rect 1790 -9480 1800 -9370
rect 1880 -9376 1890 -9318
rect 1990 -9376 2000 -9318
rect 2480 -9376 2490 -9318
rect 2590 -9376 2600 -9318
rect 2900 -9320 2910 -9220
rect 2970 -9320 2980 -9220
rect 2290 -9470 2300 -9380
rect 2360 -9470 2370 -9380
rect 2900 -9480 2910 -9370
rect 2970 -9480 2980 -9370
rect 3080 -9376 3090 -9318
rect 3190 -9376 3200 -9318
rect 3490 -9320 3500 -9220
rect 3560 -9320 3570 -9220
rect 3490 -9470 3500 -9370
rect 3560 -9470 3570 -9370
rect 3680 -9376 3690 -9318
rect 3790 -9376 3800 -9318
rect 1840 -9550 2090 -9480
rect 2190 -9550 2200 -9480
rect 2400 -9540 2690 -9480
rect 2790 -9540 2800 -9480
rect 3010 -9540 3290 -9480
rect 3390 -9500 3400 -9480
rect 3830 -9500 3880 -9220
rect 5950 -9320 5960 -9220
rect 6020 -9320 6030 -9220
rect 5210 -9380 5220 -9320
rect 5320 -9380 5330 -9320
rect 5960 -9480 6030 -9320
rect 3390 -9540 3880 -9500
rect 5410 -9540 5420 -9480
rect 5520 -9540 5530 -9480
rect 3290 -9560 3880 -9540
rect 1620 -9600 4230 -9590
rect 1620 -9640 1670 -9600
rect 4180 -9640 4230 -9600
rect 1620 -9650 4230 -9640
rect 1620 -9820 4010 -9810
rect 1620 -9860 1670 -9820
rect 3960 -9860 4010 -9820
rect 1620 -9870 4010 -9860
rect 1620 -10340 1680 -9870
rect 1960 -9960 1970 -9900
rect 2070 -9960 2080 -9900
rect 1870 -10340 1960 -10000
rect 2250 -10030 2260 -9960
rect 2390 -10030 2400 -9960
rect 2060 -10160 2070 -10030
rect 2130 -10160 2140 -10030
rect 2190 -10340 2270 -10060
rect 2370 -10250 2380 -10150
rect 2440 -10250 2450 -10150
rect 3950 -10340 4010 -9870
rect 1620 -10350 4010 -10340
rect 1620 -10390 1670 -10350
rect 3960 -10390 4010 -10350
rect 1620 -10430 4010 -10390
rect 4170 -10340 4230 -9650
rect 5010 -9680 5020 -9580
rect 5120 -9680 5710 -9580
rect 4400 -9840 4410 -9770
rect 4520 -9840 4530 -9770
rect 4560 -9840 4570 -9770
rect 4680 -9840 4690 -9770
rect 4720 -9840 4730 -9770
rect 4840 -9840 4850 -9770
rect 4350 -10150 4410 -9880
rect 4500 -10050 4510 -9950
rect 4580 -10050 4590 -9950
rect 4670 -10150 4730 -9880
rect 5330 -9940 5390 -9680
rect 5480 -9890 5490 -9790
rect 5550 -9890 5560 -9790
rect 5650 -9930 5710 -9680
rect 5800 -9890 5810 -9790
rect 5870 -9890 5880 -9790
rect 4820 -10050 4830 -9950
rect 4900 -10050 4910 -9950
rect 5370 -10050 5530 -9980
rect 5680 -10050 5920 -9980
rect 4350 -10250 5020 -10150
rect 5120 -10250 5130 -10150
rect 6060 -10340 6120 -8950
rect 4170 -10350 6120 -10340
rect 4170 -10390 4220 -10350
rect 6050 -10390 6120 -10350
rect 4170 -10400 6120 -10390
rect 1150 -10630 6130 -10430
rect 6160 -10630 6560 -8950
<< via1 >>
rect 1700 -3600 1770 -3500
rect 5950 -3600 6020 -3500
rect 2360 -3660 2460 -3600
rect 5220 -3660 5320 -3600
rect 2360 -4140 2460 -4080
rect 5220 -4140 5320 -4080
rect 2960 -4300 3060 -4240
rect 4460 -4300 4560 -4240
rect 1700 -4400 1770 -4300
rect 5960 -4400 6020 -4300
rect 2360 -4460 2460 -4400
rect 5220 -4460 5320 -4400
rect 2960 -4620 3060 -4560
rect 4460 -4620 4560 -4560
rect 2960 -4740 3060 -4680
rect 4460 -4740 4560 -4680
rect 2360 -4900 2460 -4840
rect 5220 -4900 5320 -4840
rect 1700 -5000 1770 -4900
rect 5960 -5000 6020 -4900
rect 2960 -5060 3060 -5000
rect 4460 -5060 4560 -5000
rect 2360 -5220 2460 -5160
rect 5220 -5220 5320 -5160
rect 2360 -5680 2460 -5620
rect 5220 -5680 5320 -5620
rect 1700 -5780 1770 -5680
rect 5950 -5780 6020 -5680
rect 1700 -6060 1770 -5960
rect 5950 -6060 6020 -5960
rect 2360 -6120 2460 -6060
rect 5220 -6120 5320 -6060
rect 2360 -6600 2460 -6540
rect 5220 -6600 5320 -6540
rect 2960 -6760 3060 -6700
rect 4460 -6760 4560 -6700
rect 1700 -6860 1770 -6760
rect 5960 -6860 6020 -6760
rect 2360 -6920 2460 -6860
rect 5220 -6920 5320 -6860
rect 2960 -7080 3060 -7020
rect 4460 -7080 4560 -7020
rect 2960 -7200 3060 -7140
rect 4460 -7200 4560 -7140
rect 2290 -7360 2390 -7300
rect 5220 -7360 5320 -7300
rect 1700 -7460 1770 -7360
rect 5960 -7460 6020 -7360
rect 2960 -7520 3060 -7460
rect 4460 -7520 4560 -7460
rect 2290 -7680 2390 -7620
rect 5220 -7680 5320 -7620
rect 1890 -7960 1990 -7880
rect 2490 -7960 2590 -7860
rect 3090 -7960 3190 -7860
rect 1890 -7980 1990 -7960
rect 2290 -8140 2390 -8080
rect 5220 -8140 5320 -8080
rect 1700 -8240 1770 -8140
rect 5950 -8240 6020 -8140
rect 1890 -8420 1990 -8360
rect 2490 -8420 2590 -8360
rect 3090 -8420 3190 -8360
rect 5220 -8420 5320 -8360
rect 1720 -8520 1790 -8420
rect 2290 -8510 2350 -8420
rect 2900 -8520 2960 -8420
rect 3500 -8520 3560 -8420
rect 5950 -8520 6020 -8420
rect 1890 -8580 1990 -8520
rect 2490 -8580 2590 -8520
rect 3090 -8580 3190 -8520
rect 3690 -8580 3790 -8520
rect 5420 -8580 5520 -8520
rect 2090 -8850 2190 -8750
rect 2690 -8870 2790 -8770
rect 3290 -8880 3390 -8780
rect 5020 -8890 5120 -8800
rect 5020 -8900 5120 -8890
rect 1730 -9160 1790 -9050
rect 1890 -9060 1990 -9002
rect 2490 -9060 2590 -9000
rect 3090 -9060 3190 -9000
rect 3690 -9060 3790 -9000
rect 5220 -9060 5320 -9000
rect 2300 -9150 2360 -9060
rect 2910 -9160 2970 -9060
rect 3500 -9160 3560 -9060
rect 1730 -9320 1790 -9210
rect 2090 -9220 2190 -9160
rect 2690 -9220 2790 -9160
rect 3290 -9220 3390 -9160
rect 5420 -9220 5520 -9160
rect 2300 -9310 2360 -9220
rect 1730 -9480 1790 -9370
rect 1890 -9376 1990 -9318
rect 2490 -9376 2590 -9318
rect 2910 -9320 2970 -9220
rect 2300 -9470 2360 -9380
rect 2910 -9480 2970 -9370
rect 3090 -9376 3190 -9318
rect 3500 -9320 3560 -9220
rect 3500 -9470 3560 -9370
rect 3690 -9376 3790 -9318
rect 2090 -9550 2190 -9480
rect 2690 -9540 2790 -9480
rect 3290 -9540 3390 -9480
rect 5960 -9320 6020 -9220
rect 5220 -9380 5320 -9320
rect 5420 -9540 5520 -9480
rect 1970 -9960 2070 -9900
rect 2260 -10030 2390 -9960
rect 2070 -10160 2130 -10030
rect 2380 -10250 2440 -10150
rect 5020 -9680 5120 -9580
rect 4410 -9840 4520 -9770
rect 4570 -9840 4680 -9770
rect 4730 -9840 4840 -9770
rect 4510 -10050 4580 -9950
rect 5490 -9890 5550 -9790
rect 5810 -9890 5870 -9790
rect 4830 -10050 4900 -9950
rect 5530 -10050 5680 -9980
rect 5020 -10250 5120 -10150
<< metal2 >>
rect 1090 -4300 1190 -3170
rect 1090 -4900 1190 -4400
rect 1090 -5960 1190 -5000
rect 1090 -8140 1190 -6060
rect 1090 -9110 1190 -8240
rect 1090 -10630 1190 -9210
rect 1290 -3500 1390 -3170
rect 1290 -5680 1390 -3600
rect 1290 -6760 1390 -5780
rect 1290 -7360 1390 -6860
rect 1290 -8910 1390 -7460
rect 1290 -10630 1390 -9010
rect 1490 -8710 1590 -3170
rect 1700 -3500 1770 -3490
rect 1700 -3610 1770 -3600
rect 2360 -3600 2460 -3430
rect 2360 -3790 2460 -3660
rect 2360 -4080 2460 -3890
rect 5220 -3600 5320 -3440
rect 5950 -3500 6020 -3490
rect 5950 -3610 6020 -3600
rect 1700 -4300 1770 -4290
rect 1700 -4410 1770 -4400
rect 2360 -4400 2460 -4140
rect 2360 -4620 2460 -4460
rect 2960 -3990 3060 -3980
rect 2960 -4240 3060 -4090
rect 2960 -4560 3060 -4300
rect 2960 -4630 3060 -4620
rect 4460 -3990 4560 -3980
rect 4460 -4240 4560 -4090
rect 4460 -4560 4560 -4300
rect 4460 -4630 4560 -4620
rect 5220 -4080 5320 -3660
rect 5220 -4400 5320 -4140
rect 5960 -4300 6020 -4290
rect 5960 -4410 6020 -4400
rect 2960 -4680 3060 -4670
rect 2360 -4840 2460 -4680
rect 1700 -4900 1770 -4890
rect 1700 -5010 1770 -5000
rect 2360 -5160 2460 -4900
rect 2360 -5400 2460 -5220
rect 2960 -5000 3060 -4740
rect 2960 -5200 3060 -5060
rect 2960 -5310 3060 -5300
rect 4460 -4680 4560 -4670
rect 4460 -5000 4560 -4740
rect 4460 -5200 4560 -5060
rect 4460 -5310 4560 -5300
rect 5220 -4840 5320 -4460
rect 5220 -5160 5320 -4900
rect 5960 -4900 6020 -4890
rect 5960 -5010 6020 -5000
rect 2360 -5620 2460 -5500
rect 1700 -5680 1770 -5670
rect 1700 -5790 1770 -5780
rect 2360 -5840 2460 -5680
rect 5220 -5620 5320 -5220
rect 1700 -5960 1770 -5950
rect 1700 -6070 1770 -6060
rect 2360 -6060 2460 -5900
rect 2360 -6250 2460 -6120
rect 5220 -6060 5320 -5680
rect 5950 -5680 6020 -5670
rect 5950 -5790 6020 -5780
rect 5950 -5960 6020 -5950
rect 5950 -6070 6020 -6060
rect 2460 -6310 2470 -6250
rect 2360 -6540 2460 -6350
rect 1700 -6760 1770 -6750
rect 1700 -6870 1770 -6860
rect 2360 -6860 2460 -6600
rect 2360 -7080 2460 -6920
rect 2960 -6450 3060 -6440
rect 2960 -6700 3060 -6550
rect 2960 -7020 3060 -6760
rect 2960 -7090 3060 -7080
rect 4460 -6450 4560 -6440
rect 4460 -6700 4560 -6550
rect 4460 -7020 4560 -6760
rect 4460 -7090 4560 -7080
rect 5220 -6540 5320 -6120
rect 5220 -6860 5320 -6600
rect 5960 -6760 6020 -6750
rect 5960 -6870 6020 -6860
rect 2960 -7140 3060 -7130
rect 2290 -7300 2390 -7140
rect 1700 -7360 1770 -7350
rect 1700 -7470 1770 -7460
rect 2290 -7620 2390 -7360
rect 2290 -7860 2390 -7680
rect 2960 -7460 3060 -7200
rect 2960 -7660 3060 -7520
rect 2960 -7770 3060 -7760
rect 4460 -7140 4560 -7130
rect 4460 -7460 4560 -7200
rect 4460 -7660 4560 -7520
rect 4460 -7770 4560 -7760
rect 5220 -7300 5320 -6920
rect 5220 -7620 5320 -7360
rect 5960 -7360 6020 -7350
rect 5960 -7470 6020 -7460
rect 1890 -7880 1990 -7870
rect 1700 -8140 1770 -8130
rect 1700 -8250 1770 -8240
rect 1890 -8360 1990 -7980
rect 2290 -8080 2390 -7960
rect 2290 -8300 2390 -8140
rect 2490 -7860 2590 -7850
rect 1490 -10630 1590 -8810
rect 1690 -8420 1790 -8400
rect 1690 -8520 1720 -8420
rect 2490 -8360 2590 -7960
rect 1890 -8430 1990 -8420
rect 2290 -8420 2390 -8390
rect 1690 -8710 1790 -8520
rect 1690 -9050 1790 -8810
rect 1690 -9160 1730 -9050
rect 1690 -9210 1790 -9160
rect 1690 -9320 1730 -9210
rect 1690 -9370 1790 -9320
rect 1690 -9480 1730 -9370
rect 1690 -9490 1790 -9480
rect 1890 -8520 1990 -8500
rect 1890 -8910 1990 -8580
rect 2350 -8510 2390 -8420
rect 3090 -7860 3190 -7850
rect 3090 -8360 3190 -7960
rect 2900 -8420 2960 -8410
rect 3690 -7860 3790 -7850
rect 2490 -8430 2590 -8420
rect 1890 -9318 1990 -9060
rect 1890 -9540 1990 -9376
rect 2090 -8750 2190 -8620
rect 2090 -9160 2190 -8850
rect 2090 -9480 2190 -9220
rect 2290 -8910 2390 -8510
rect 2290 -9060 2390 -9010
rect 2290 -9150 2300 -9060
rect 2360 -9150 2390 -9060
rect 2290 -9220 2390 -9150
rect 2290 -9310 2300 -9220
rect 2360 -9310 2390 -9220
rect 2290 -9380 2390 -9310
rect 2290 -9470 2300 -9380
rect 2360 -9470 2390 -9380
rect 2290 -9540 2390 -9470
rect 2490 -8520 2590 -8510
rect 2490 -9000 2590 -8580
rect 2890 -8520 2900 -8420
rect 2960 -8520 2990 -8420
rect 3090 -8430 3190 -8420
rect 3490 -8420 3590 -8370
rect 2490 -9110 2590 -9060
rect 2490 -9318 2590 -9210
rect 2490 -9540 2590 -9376
rect 2690 -8770 2790 -8620
rect 2690 -9160 2790 -8870
rect 2690 -9480 2790 -9220
rect 2890 -8720 2990 -8520
rect 2890 -9060 2990 -8810
rect 2890 -9160 2910 -9060
rect 2970 -9160 2990 -9060
rect 2890 -9220 2990 -9160
rect 2890 -9320 2910 -9220
rect 2970 -9320 2990 -9220
rect 2890 -9370 2990 -9320
rect 2890 -9480 2910 -9370
rect 2970 -9480 2990 -9370
rect 2890 -9540 2990 -9480
rect 3090 -8520 3190 -8510
rect 3090 -9000 3190 -8580
rect 3490 -8520 3500 -8420
rect 3560 -8520 3590 -8420
rect 3090 -9318 3190 -9060
rect 2690 -9550 2790 -9540
rect 3090 -9550 3190 -9376
rect 3290 -8780 3390 -8620
rect 3290 -9160 3390 -8880
rect 3290 -9480 3390 -9220
rect 3290 -9550 3390 -9540
rect 3490 -9060 3590 -8520
rect 3490 -9160 3500 -9060
rect 3560 -9160 3590 -9060
rect 3490 -9220 3590 -9160
rect 3490 -9320 3500 -9220
rect 3560 -9320 3590 -9220
rect 3490 -9370 3590 -9320
rect 3490 -9470 3500 -9370
rect 3560 -9470 3590 -9370
rect 3490 -9550 3590 -9470
rect 3690 -8520 3790 -7960
rect 3690 -9000 3790 -8580
rect 5220 -8080 5320 -7680
rect 5220 -8360 5320 -8140
rect 5950 -8140 6020 -8130
rect 5950 -8250 6020 -8240
rect 3690 -9318 3790 -9060
rect 3690 -9540 3790 -9376
rect 5020 -8800 5120 -8790
rect 2090 -9560 2190 -9550
rect 3090 -9660 3190 -9650
rect 3490 -9660 3590 -9650
rect 5020 -9580 5120 -8900
rect 5220 -9000 5320 -8420
rect 5220 -9320 5320 -9060
rect 5220 -9540 5320 -9380
rect 5420 -8520 5520 -8360
rect 5950 -8420 6020 -8410
rect 5950 -8530 6020 -8520
rect 5420 -8910 5520 -8580
rect 5420 -9160 5520 -9010
rect 6130 -8720 6230 -3170
rect 5420 -9480 5520 -9220
rect 5960 -9220 6020 -9210
rect 5960 -9330 6020 -9320
rect 5420 -9550 5520 -9540
rect 1970 -9750 2070 -9740
rect 4410 -9770 4520 -9760
rect 4410 -9850 4520 -9840
rect 4570 -9770 4680 -9760
rect 4570 -9850 4680 -9840
rect 4730 -9770 4840 -9760
rect 4730 -9850 4840 -9840
rect 1970 -9900 2070 -9850
rect 4510 -9950 4580 -9940
rect 1970 -9970 2070 -9960
rect 2260 -9960 2390 -9950
rect 2070 -10030 2130 -10020
rect 2260 -10040 2390 -10030
rect 4510 -10060 4580 -10050
rect 4830 -9950 4900 -9940
rect 4830 -10060 4900 -10050
rect 2070 -10170 2130 -10160
rect 2380 -10150 2440 -10140
rect 2380 -10260 2440 -10250
rect 5020 -10150 5120 -9680
rect 5490 -9790 5550 -9780
rect 5810 -9790 5870 -9780
rect 5020 -10260 5120 -10250
rect 5220 -9890 5490 -9790
rect 5550 -9890 5810 -9790
rect 5870 -9890 5890 -9790
rect 5220 -10150 5320 -9890
rect 5490 -9900 5550 -9890
rect 5810 -9900 5870 -9890
rect 5530 -9980 5680 -9970
rect 5530 -10060 5680 -10050
rect 5220 -10260 5320 -10250
rect 6130 -10630 6230 -8810
rect 6330 -3500 6430 -3170
rect 6330 -4900 6430 -3600
rect 6330 -5960 6430 -5000
rect 6330 -7360 6430 -6060
rect 6330 -9550 6430 -7460
rect 6330 -10630 6430 -9650
rect 6530 -4300 6630 -3170
rect 6530 -5680 6630 -4400
rect 6530 -6760 6630 -5780
rect 6530 -7860 6630 -6860
rect 6530 -8140 6630 -7960
rect 6530 -10630 6630 -8240
rect 6730 -9750 6830 -3170
rect 6730 -10630 6830 -9850
rect 6930 -9220 7030 -3170
rect 6930 -9950 7030 -9320
rect 6930 -10630 7030 -10050
rect 7130 -8420 7230 -3170
rect 7130 -10150 7230 -8520
rect 7130 -10630 7230 -10250
<< via2 >>
rect 1090 -4400 1190 -4300
rect 1090 -5000 1190 -4900
rect 1090 -6060 1190 -5960
rect 1090 -8240 1190 -8140
rect 1090 -9210 1190 -9110
rect 1290 -3600 1390 -3500
rect 1290 -5780 1390 -5680
rect 1290 -6860 1390 -6760
rect 1290 -7460 1390 -7360
rect 1290 -9010 1390 -8910
rect 1700 -3600 1770 -3500
rect 2360 -3890 2460 -3790
rect 5950 -3600 6020 -3500
rect 1700 -4400 1770 -4300
rect 2960 -4090 3060 -3990
rect 4460 -4090 4560 -3990
rect 5960 -4400 6020 -4300
rect 1700 -5000 1770 -4900
rect 2960 -5300 3060 -5200
rect 4460 -5300 4560 -5200
rect 5960 -5000 6020 -4900
rect 2360 -5500 2460 -5400
rect 1700 -5780 1770 -5680
rect 1700 -6060 1770 -5960
rect 5950 -5780 6020 -5680
rect 5950 -6060 6020 -5960
rect 2360 -6350 2460 -6250
rect 1700 -6860 1770 -6760
rect 2960 -6550 3060 -6450
rect 4460 -6550 4560 -6450
rect 5960 -6860 6020 -6760
rect 1700 -7460 1770 -7360
rect 2960 -7760 3060 -7660
rect 4460 -7760 4560 -7660
rect 5960 -7460 6020 -7360
rect 1700 -8240 1770 -8140
rect 2290 -7960 2390 -7860
rect 1490 -8810 1590 -8710
rect 1690 -8810 1790 -8710
rect 3690 -7960 3790 -7860
rect 1890 -9002 1990 -8910
rect 1890 -9010 1990 -9002
rect 2290 -9010 2390 -8910
rect 2490 -9210 2590 -9110
rect 2890 -8810 2990 -8720
rect 5950 -8240 6020 -8140
rect 3090 -9650 3190 -9550
rect 3490 -9650 3590 -9550
rect 5950 -8520 6020 -8420
rect 5420 -9010 5520 -8910
rect 6130 -8810 6230 -8720
rect 5960 -9320 6020 -9220
rect 1970 -9850 2070 -9750
rect 4410 -9840 4520 -9770
rect 4570 -9840 4680 -9770
rect 4730 -9840 4840 -9770
rect 2070 -10160 2130 -10030
rect 2260 -10030 2390 -9960
rect 4510 -10050 4580 -9950
rect 4830 -10050 4900 -9950
rect 2380 -10250 2440 -10150
rect 5530 -10050 5680 -9980
rect 5220 -10250 5320 -10150
rect 6330 -3600 6430 -3500
rect 6330 -5000 6430 -4900
rect 6330 -6060 6430 -5960
rect 6330 -7460 6430 -7360
rect 6330 -9650 6430 -9550
rect 6530 -4400 6630 -4300
rect 6530 -5780 6630 -5680
rect 6530 -6860 6630 -6760
rect 6530 -7960 6630 -7860
rect 6530 -8240 6630 -8140
rect 6730 -9850 6830 -9750
rect 6930 -9320 7030 -9220
rect 6930 -10050 7030 -9950
rect 7130 -8520 7230 -8420
rect 7130 -10250 7230 -10150
<< metal3 >>
rect 1280 -3500 1400 -3495
rect 1690 -3500 1780 -3495
rect 1280 -3600 1290 -3500
rect 1390 -3600 1700 -3500
rect 1770 -3600 1780 -3500
rect 1280 -3605 1400 -3600
rect 1690 -3605 1780 -3600
rect 5940 -3500 6030 -3495
rect 6320 -3500 6440 -3495
rect 5940 -3600 5950 -3500
rect 6020 -3600 6330 -3500
rect 6430 -3600 6440 -3500
rect 5940 -3605 6030 -3600
rect 6320 -3605 6440 -3600
rect 2350 -3790 2470 -3785
rect 990 -3890 2360 -3790
rect 2460 -3890 3820 -3790
rect 2350 -3895 2470 -3890
rect 2950 -3990 3070 -3985
rect 4450 -3990 4570 -3985
rect 2950 -4090 2960 -3990
rect 3060 -4090 4460 -3990
rect 4560 -4090 4570 -3990
rect 2950 -4095 3070 -4090
rect 4450 -4095 4570 -4090
rect 1080 -4300 1200 -4295
rect 1690 -4300 1780 -4295
rect 1080 -4400 1090 -4300
rect 1190 -4400 1700 -4300
rect 1770 -4400 1780 -4300
rect 1080 -4405 1200 -4400
rect 1690 -4405 1780 -4400
rect 5950 -4300 6030 -4295
rect 6520 -4300 6640 -4295
rect 5950 -4400 5960 -4300
rect 6020 -4400 6530 -4300
rect 6630 -4400 6640 -4300
rect 5950 -4405 6030 -4400
rect 6520 -4405 6640 -4400
rect 1080 -4900 1200 -4895
rect 1690 -4900 1780 -4895
rect 1080 -5000 1090 -4900
rect 1190 -5000 1700 -4900
rect 1770 -5000 1780 -4900
rect 1080 -5005 1200 -5000
rect 1690 -5005 1780 -5000
rect 5950 -4900 6030 -4895
rect 6320 -4900 6440 -4895
rect 5950 -5000 5960 -4900
rect 6020 -5000 6330 -4900
rect 6430 -5000 6440 -4900
rect 5950 -5005 6030 -5000
rect 6320 -5005 6440 -5000
rect 2950 -5200 3070 -5195
rect 4450 -5200 4570 -5195
rect 2950 -5300 2960 -5200
rect 3060 -5300 4460 -5200
rect 4560 -5300 4570 -5200
rect 2950 -5305 3070 -5300
rect 4450 -5305 4570 -5300
rect 2350 -5400 2470 -5395
rect 990 -5500 2360 -5400
rect 2460 -5500 3820 -5400
rect 2350 -5505 2470 -5500
rect 1280 -5680 1400 -5675
rect 1690 -5680 1780 -5675
rect 1280 -5780 1290 -5680
rect 1390 -5780 1700 -5680
rect 1770 -5780 1780 -5680
rect 1280 -5785 1400 -5780
rect 1690 -5785 1780 -5780
rect 5940 -5680 6030 -5675
rect 6520 -5680 6640 -5675
rect 5940 -5780 5950 -5680
rect 6020 -5780 6530 -5680
rect 6630 -5780 6640 -5680
rect 5940 -5785 6030 -5780
rect 6520 -5785 6640 -5780
rect 1080 -5960 1200 -5955
rect 1690 -5960 1780 -5955
rect 1080 -6060 1090 -5960
rect 1190 -6060 1700 -5960
rect 1770 -6060 1780 -5960
rect 1080 -6065 1200 -6060
rect 1690 -6065 1780 -6060
rect 5940 -5960 6030 -5955
rect 6320 -5960 6440 -5955
rect 5940 -6060 5950 -5960
rect 6020 -6060 6330 -5960
rect 6430 -6060 6440 -5960
rect 5940 -6065 6030 -6060
rect 6320 -6065 6440 -6060
rect 2350 -6250 2470 -6245
rect 990 -6350 2360 -6250
rect 2460 -6350 3820 -6250
rect 2350 -6355 2470 -6350
rect 2950 -6450 3070 -6445
rect 4450 -6450 4570 -6445
rect 2950 -6550 2960 -6450
rect 3060 -6550 4460 -6450
rect 4560 -6550 4570 -6450
rect 2950 -6555 3070 -6550
rect 4450 -6555 4570 -6550
rect 1280 -6760 1400 -6755
rect 1690 -6760 1780 -6755
rect 1280 -6860 1290 -6760
rect 1390 -6860 1700 -6760
rect 1770 -6860 1780 -6760
rect 1280 -6865 1400 -6860
rect 1690 -6865 1780 -6860
rect 5950 -6760 6030 -6755
rect 6520 -6760 6640 -6755
rect 5950 -6860 5960 -6760
rect 6020 -6860 6530 -6760
rect 6630 -6860 6640 -6760
rect 5950 -6865 6030 -6860
rect 6520 -6865 6640 -6860
rect 1280 -7360 1400 -7355
rect 1690 -7360 1780 -7355
rect 1280 -7460 1290 -7360
rect 1390 -7460 1700 -7360
rect 1770 -7460 1780 -7360
rect 1280 -7465 1400 -7460
rect 1690 -7465 1780 -7460
rect 5950 -7360 6030 -7355
rect 6320 -7360 6440 -7355
rect 5950 -7460 5960 -7360
rect 6020 -7460 6330 -7360
rect 6430 -7460 6440 -7360
rect 5950 -7465 6030 -7460
rect 6320 -7465 6440 -7460
rect 2950 -7660 3070 -7655
rect 4450 -7660 4570 -7655
rect 2950 -7760 2960 -7660
rect 3060 -7760 4460 -7660
rect 4560 -7760 4570 -7660
rect 2950 -7765 3070 -7760
rect 4450 -7765 4570 -7760
rect 2280 -7860 2400 -7855
rect 3680 -7860 3800 -7855
rect 6520 -7860 6640 -7855
rect 990 -7960 2290 -7860
rect 2390 -7960 2710 -7860
rect 2960 -7960 3690 -7860
rect 3790 -7960 6530 -7860
rect 6630 -7960 6640 -7860
rect 2280 -7965 2400 -7960
rect 3680 -7965 3800 -7960
rect 6520 -7965 6640 -7960
rect 1080 -8140 1200 -8135
rect 1690 -8140 1780 -8135
rect 1080 -8240 1090 -8140
rect 1190 -8240 1700 -8140
rect 1770 -8240 1780 -8140
rect 1080 -8245 1200 -8240
rect 1690 -8245 1780 -8240
rect 5940 -8140 6030 -8135
rect 6520 -8140 6640 -8135
rect 5940 -8240 5950 -8140
rect 6020 -8240 6530 -8140
rect 6630 -8240 6640 -8140
rect 5940 -8245 6030 -8240
rect 6520 -8245 6640 -8240
rect 5940 -8420 6030 -8415
rect 7120 -8420 7240 -8415
rect 5940 -8520 5950 -8420
rect 6020 -8520 7130 -8420
rect 7230 -8520 7240 -8420
rect 5940 -8525 6030 -8520
rect 7120 -8525 7240 -8520
rect 1480 -8710 1600 -8705
rect 1680 -8710 1800 -8705
rect 1480 -8810 1490 -8710
rect 1590 -8810 1690 -8710
rect 1790 -8810 1800 -8710
rect 1480 -8815 1600 -8810
rect 1680 -8815 1800 -8810
rect 2880 -8720 3000 -8715
rect 6120 -8720 6240 -8715
rect 2880 -8810 2890 -8720
rect 2990 -8810 6130 -8720
rect 6230 -8810 6240 -8720
rect 2880 -8815 3000 -8810
rect 6120 -8815 6240 -8810
rect 1280 -8910 1400 -8905
rect 1880 -8910 2000 -8905
rect 2280 -8910 2400 -8905
rect 5410 -8910 5530 -8905
rect 1280 -9010 1290 -8910
rect 1390 -9010 1890 -8910
rect 1990 -9010 2290 -8910
rect 2390 -9010 2400 -8910
rect 3910 -9010 5420 -8910
rect 5520 -9010 7330 -8910
rect 1280 -9015 1400 -9010
rect 1880 -9015 2000 -9010
rect 2280 -9015 2400 -9010
rect 5410 -9015 5530 -9010
rect 1080 -9110 1200 -9105
rect 2480 -9110 2600 -9105
rect 1080 -9210 1090 -9110
rect 1190 -9210 2490 -9110
rect 2590 -9210 2600 -9110
rect 1080 -9215 1200 -9210
rect 2480 -9215 2600 -9210
rect 5950 -9220 6030 -9215
rect 6920 -9220 7040 -9215
rect 5950 -9320 5960 -9220
rect 6020 -9320 6930 -9220
rect 7030 -9320 7040 -9220
rect 5950 -9325 6030 -9320
rect 6920 -9325 7040 -9320
rect 3080 -9550 3200 -9545
rect 3480 -9550 3600 -9545
rect 6320 -9550 6440 -9545
rect 3080 -9650 3090 -9550
rect 3190 -9650 3490 -9550
rect 3590 -9650 6330 -9550
rect 6430 -9650 6440 -9550
rect 3080 -9655 3200 -9650
rect 3480 -9655 3600 -9650
rect 6320 -9655 6440 -9650
rect 1960 -9750 2080 -9745
rect 6720 -9750 6840 -9745
rect 1930 -9850 1970 -9750
rect 2070 -9770 6730 -9750
rect 2070 -9840 4410 -9770
rect 4520 -9840 4570 -9770
rect 4680 -9840 4730 -9770
rect 4840 -9840 6730 -9770
rect 2070 -9850 6730 -9840
rect 6830 -9850 6840 -9750
rect 1960 -9855 2080 -9850
rect 6720 -9855 6840 -9850
rect 4500 -9950 4590 -9945
rect 2070 -9960 4410 -9950
rect 4500 -9960 4510 -9950
rect 2070 -10025 2260 -9960
rect 2060 -10030 2260 -10025
rect 2390 -10030 4510 -9960
rect 2060 -10160 2070 -10030
rect 2130 -10050 4510 -10030
rect 4580 -9960 4590 -9950
rect 4820 -9950 4910 -9945
rect 6920 -9950 7040 -9945
rect 4820 -9960 4830 -9950
rect 4580 -10050 4830 -9960
rect 4900 -9980 6930 -9950
rect 4900 -10050 5530 -9980
rect 5680 -10050 6930 -9980
rect 7030 -10050 7040 -9950
rect 2130 -10160 2140 -10050
rect 4500 -10055 4590 -10050
rect 4820 -10055 4910 -10050
rect 5520 -10055 5690 -10050
rect 6920 -10055 7040 -10050
rect 2060 -10165 2140 -10160
rect 2370 -10150 2450 -10145
rect 5210 -10150 5330 -10145
rect 7120 -10150 7240 -10145
rect 2370 -10250 2380 -10150
rect 2440 -10250 5220 -10150
rect 5320 -10250 7130 -10150
rect 7230 -10250 7240 -10150
rect 2370 -10255 2450 -10250
rect 5210 -10255 5330 -10250
rect 7120 -10255 7240 -10250
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM1
timestamp 1736329344
transform 0 -1 2779 1 0 -5732
box -108 -1057 108 1057
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM2
timestamp 1736329344
transform 0 -1 2774 1 0 -4948
box -332 -1102 332 1064
use sky130_fd_pr__nfet_g5v0d10v5_SMV9TY  XM3
timestamp 1736329706
transform 0 -1 3667 1 0 -8472
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_KNBJVF  XM4
timestamp 1736363543
transform 0 -1 3664 1 0 -9268
box -332 -202 332 164
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM5
timestamp 1736329344
transform 0 -1 2779 1 0 -3552
box -108 -1057 108 1057
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM6
timestamp 1736329344
transform 0 -1 2774 -1 0 -4348
box -332 -1102 332 1064
use sky130_fd_pr__nfet_g5v0d10v5_SMV9TY  XM7
timestamp 1736329706
transform 0 -1 3067 1 0 -8472
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_KNBJVF  XM8
timestamp 1736363543
transform 0 -1 3074 1 0 -9268
box -332 -202 332 164
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM9
timestamp 1736329344
transform 0 -1 2779 -1 0 -8192
box -108 -1057 108 1057
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM10
timestamp 1736329344
transform 0 -1 2774 1 0 -7408
box -332 -1102 332 1064
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM11
timestamp 1736329344
transform 0 1 4946 -1 0 -4348
box -332 -1102 332 1064
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM12
timestamp 1736329344
transform 0 1 4941 -1 0 -3552
box -108 -1057 108 1057
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM13
timestamp 1736329344
transform 0 -1 2779 1 0 -6012
box -108 -1057 108 1057
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM14
timestamp 1736329344
transform 0 -1 2774 1 0 -6808
box -332 -1102 332 1064
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM15
timestamp 1736329344
transform 0 1 4946 -1 0 -4948
box -332 -1102 332 1064
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM16
timestamp 1736329344
transform 0 1 4941 -1 0 -5732
box -108 -1057 108 1057
use sky130_fd_pr__nfet_g5v0d10v5_SMV9TY  XM17
timestamp 1736329706
transform 0 -1 2457 -1 0 -8472
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_KNBJVF  XM18
timestamp 1736363543
transform 0 -1 2464 1 0 -9268
box -332 -202 332 164
use sky130_fd_pr__nfet_g5v0d10v5_SMV9TY  XM19
timestamp 1736329706
transform 0 -1 1897 1 0 -8472
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_KNBJVF  XM20
timestamp 1736363543
transform 0 -1 1904 -1 0 -9268
box -332 -202 332 164
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM21
timestamp 1736329344
transform 0 1 4946 -1 0 -6808
box -332 -1102 332 1064
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM22
timestamp 1736329344
transform 0 1 4941 -1 0 -6012
box -108 -1057 108 1057
use sky130_fd_pr__pfet_g5v0d10v5_PE8P5C  XM23
timestamp 1736329344
transform 0 1 4946 1 0 -7408
box -332 -1102 332 1064
use sky130_fd_pr__nfet_g5v0d10v5_H5TWCS  XM24
timestamp 1736329344
transform 0 1 4941 -1 0 -8192
box -108 -1057 108 1057
use sky130_fd_pr__pfet_g5v0d10v5_K2M7HA  XM25
timestamp 1736363715
transform 0 1 4946 -1 0 -9268
box -332 -1102 332 1064
use sky130_fd_pr__nfet_g5v0d10v5_Y8DDSH  XM26
timestamp 1736339096
transform 0 -1 4941 1 0 -8472
box -108 -1057 108 1057
use sky130_fd_pr__nfet_g5v0d10v5_Z6HFXJ  XM27
timestamp 1736338749
transform 1 0 2328 0 1 -10133
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_K8GQEA  XM28
timestamp 1736363663
transform -1 0 5602 0 -1 -9876
box -332 -202 332 164
use sky130_fd_pr__nfet_g5v0d10v5_Z6HFXJ  XM29
timestamp 1736338749
transform -1 0 2018 0 1 -10063
box -108 -157 108 157
use sky130_fd_pr__pfet_g5v0d10v5_K8GQEA  XM30
timestamp 1736363663
transform -1 0 4622 0 1 -9938
box -332 -202 332 164
<< labels >>
flabel metal3 990 -3890 1090 -3790 0 FreeSans 160 0 0 0 mux_inA
port 10 nsew
flabel metal3 990 -5500 1090 -5400 0 FreeSans 160 0 0 0 mux_inB
port 16 nsew
flabel metal3 990 -6350 1090 -6250 0 FreeSans 160 0 0 0 mux_inC
port 17 nsew
flabel metal3 990 -7960 1090 -7860 0 FreeSans 160 0 0 0 mux_inD
port 18 nsew
flabel metal3 7230 -9010 7330 -8910 0 FreeSans 160 0 0 0 mux_out
port 30 nsew
flabel metal1 1150 -3270 1250 -3170 0 FreeSans 160 0 0 0 vssa
port 45 nsew
flabel metal1 6460 -3270 6560 -3170 0 FreeSans 160 0 0 0 vdda
port 44 nsew
flabel metal2 1490 -10630 1590 -10530 0 FreeSans 160 0 0 0 sel1
port 7 nsew
flabel metal2 6130 -10630 6230 -10530 0 FreeSans 160 0 0 0 sel0
port 5 nsew
flabel metal2 6730 -10630 6830 -10530 0 FreeSans 160 0 0 0 ena
port 50 nsew
<< end >>
