magic
tech sky130A
magscale 1 2
timestamp 1736253881
<< metal3 >>
rect -1886 3012 1886 3040
rect -1886 -3012 1802 3012
rect 1866 -3012 1886 3012
rect -1886 -3040 1886 -3012
<< via3 >>
rect 1802 -3012 1866 3012
<< mimcap >>
rect -1846 2960 1554 3000
rect -1846 -2960 -1806 2960
rect 1514 -2960 1554 2960
rect -1846 -3000 1554 -2960
<< mimcapcontact >>
rect -1806 -2960 1514 2960
<< metal4 >>
rect 1786 3012 1882 3028
rect -1807 2960 1515 2961
rect -1807 -2960 -1806 2960
rect 1514 -2960 1515 2960
rect -1807 -2961 1515 -2960
rect 1786 -3012 1802 3012
rect 1866 -3012 1882 3012
rect 1786 -3028 1882 -3012
<< properties >>
string FIXED_BBOX -1886 -3040 1594 3040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 17 l 30.0 val 1.037k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
