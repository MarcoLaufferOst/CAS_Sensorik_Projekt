magic
tech sky130A
magscale 1 2
timestamp 1736177760
<< metal1 >>
rect -1190 5996 5342 5998
rect -1200 5638 -1190 5996
rect -640 5638 5342 5996
rect -1200 5634 -626 5638
rect -440 2064 -360 2080
rect -440 2060 -346 2064
rect -467 2040 -440 2058
rect -340 2042 -261 2058
rect -410 2040 -400 2042
rect -490 1960 -480 2040
rect -320 1971 -261 2042
rect 304 2040 314 2042
rect -320 1960 -310 1971
rect 252 1960 262 2040
rect 394 1960 404 2042
rect 1050 2040 1060 2042
rect 992 1960 1002 2040
rect 1140 1960 1150 2042
rect 1792 2040 1802 2042
rect 1734 1960 1744 2040
rect 1882 1960 1892 2042
rect 2538 2040 2548 2042
rect 2478 1960 2488 2040
rect 2628 1960 2638 2042
rect 3278 2040 3288 2042
rect 3222 1960 3232 2040
rect 3368 1960 3378 2042
rect 4018 2040 4028 2042
rect 3968 1960 3978 2040
rect 4108 1960 4118 2042
rect 4758 2040 4768 2042
rect 4702 1960 4712 2040
rect 4848 1960 4858 2042
rect -1186 200 5112 202
rect -1196 -40 -1186 200
rect -640 -40 5342 200
rect -1186 -442 -960 -40
rect -134 -406 -124 -206
rect 76 -406 86 -206
rect 566 -404 576 -204
rect 776 -404 786 -204
rect 1264 -402 1274 -204
rect 1476 -402 1486 -204
rect 1972 -404 1982 -204
rect 2182 -404 2192 -204
rect 2670 -402 2680 -200
rect 2884 -402 2894 -200
rect 3370 -402 3380 -200
rect 3580 -402 3590 -200
rect 4070 -404 4080 -202
rect 4282 -404 4292 -202
rect 4350 -834 4360 -202
rect 4710 -834 4720 -202
rect 4776 -402 4786 -202
rect 4986 -402 4996 -202
rect 5062 -240 5342 -40
<< via1 >>
rect -1190 5638 -640 5996
rect -400 2040 -320 2042
rect -480 1960 -320 2040
rect 314 2040 394 2042
rect 262 1960 394 2040
rect 1060 2040 1140 2042
rect 1002 1960 1140 2040
rect 1802 2040 1882 2042
rect 1744 1960 1882 2040
rect 2548 2040 2628 2042
rect 2488 1960 2628 2040
rect 3288 2040 3368 2042
rect 3232 1960 3368 2040
rect 4028 2040 4108 2042
rect 3978 1960 4108 2040
rect 4768 2040 4848 2042
rect 4712 1960 4848 2040
rect -1186 -40 -640 200
rect -124 -406 76 -206
rect 576 -404 776 -204
rect 1274 -402 1476 -204
rect 1982 -404 2182 -204
rect 2680 -402 2884 -200
rect 3380 -402 3580 -200
rect 4080 -404 4282 -202
rect 4360 -834 4710 -202
rect 4786 -402 4986 -202
<< metal2 >>
rect -1202 5996 -640 6006
rect -1202 5638 -1190 5996
rect -404 5820 -320 5998
rect -1202 5628 -640 5638
rect -403 2050 -320 5820
rect 314 2050 394 5998
rect 1060 2050 1140 5998
rect 1802 2050 1882 5998
rect 2548 2050 2628 5998
rect 3288 2050 3368 5998
rect 4028 2050 4108 5998
rect 4768 2050 4848 5998
rect -480 2042 -320 2050
rect -480 2040 -400 2042
rect -480 1950 -320 1960
rect 262 2042 394 2050
rect 262 2040 314 2042
rect 262 1950 394 1960
rect 1002 2042 1140 2050
rect 1002 2040 1060 2042
rect 1002 1950 1140 1960
rect 1744 2042 1882 2050
rect 1744 2040 1802 2042
rect 1744 1950 1882 1960
rect 2488 2042 2628 2050
rect 2488 2040 2548 2042
rect 2488 1950 2628 1960
rect 3232 2042 3368 2050
rect 3232 2040 3288 2042
rect 3232 1950 3368 1960
rect 3978 2042 4108 2050
rect 3978 2040 4028 2042
rect 3978 1950 4108 1960
rect 4712 2042 4848 2050
rect 4712 2040 4768 2042
rect 4712 1950 4848 1960
rect -1186 200 -640 210
rect -1186 -50 -640 -40
rect -484 -196 -282 200
rect 254 -194 456 202
rect 1000 -192 1198 202
rect -484 -206 78 -196
rect -484 -406 -124 -206
rect 76 -406 78 -206
rect -484 -416 78 -406
rect 254 -204 776 -194
rect 254 -404 576 -204
rect 254 -414 776 -404
rect 1000 -204 1480 -192
rect 1000 -402 1274 -204
rect 1476 -402 1480 -204
rect 1000 -412 1480 -402
rect 1738 -194 1942 202
rect 2480 -190 2680 200
rect 3224 -188 3426 202
rect 1738 -204 2182 -194
rect 1738 -404 1982 -204
rect 254 -416 774 -414
rect 1738 -416 2182 -404
rect 2480 -200 2884 -190
rect 2480 -402 2680 -200
rect 2480 -412 2884 -402
rect 3224 -200 3580 -188
rect 3224 -402 3380 -200
rect 3224 -414 3580 -402
rect 3966 -192 4166 202
rect 4708 2 4986 202
rect 3966 -202 4282 -192
rect 3966 -404 4080 -202
rect 3966 -414 4282 -404
rect 4360 -202 4710 -192
rect 4786 -202 4986 2
rect 4786 -412 4986 -402
rect 4710 -744 5342 -512
rect 4360 -844 4710 -834
<< metal4 >>
rect -961 5637 -639 5881
use dac_switch  dac_switch_0
timestamp 1736094482
transform 1 0 -1674 0 1 1446
box 742 -1446 1674 4390
use dac_switch  dac_switch_1
timestamp 1736094482
transform 1 0 -934 0 1 1448
box 742 -1446 1674 4390
use dac_switch  dac_switch_2
timestamp 1736094482
transform 1 0 -192 0 1 1448
box 742 -1446 1674 4390
use dac_switch  dac_switch_3
timestamp 1736094482
transform 1 0 550 0 1 1448
box 742 -1446 1674 4390
use dac_switch  dac_switch_4
timestamp 1736094482
transform 1 0 1292 0 1 1448
box 742 -1446 1674 4390
use dac_switch  dac_switch_5
timestamp 1736094482
transform 1 0 2034 0 1 1448
box 742 -1446 1674 4390
use dac_switch  dac_switch_6
timestamp 1736094482
transform 1 0 2776 0 1 1448
box 742 -1446 1674 4390
use dac_switch  dac_switch_7
timestamp 1736094482
transform 1 0 3518 0 1 1448
box 742 -1446 1674 4390
use R2R_20k  R2R_20k_0
timestamp 1736115234
transform 1 0 -3516 0 1 200
box 2318 -3004 8872 -400
<< labels >>
rlabel metal2 5214 -694 5346 -560 1 V_out
port 1 n
rlabel metal2 4768 5920 4848 5998 1 D7
port 2 n
rlabel metal2 -404 5920 -320 5998 1 D0
port 3 n
rlabel metal2 314 5920 394 5998 1 D1
port 4 n
rlabel metal2 4028 5920 4108 5998 1 D6
port 5 n
rlabel metal2 1060 5920 1140 5998 1 D2
port 6 n
rlabel metal2 3288 5920 3368 5998 1 D5
port 7 n
rlabel metal2 1802 5920 1882 5998 1 D3
port 8 n
rlabel metal2 2548 5920 2628 5998 1 D4
port 9 n
rlabel metal2 -1080 62 -1080 62 1 V_COM
port 11 n
rlabel metal2 -1146 5812 -1146 5812 1 V_REF
port 10 n
<< end >>
